`timescale 1ns / 1ps

module decision_tree_leaves_0(input logic [0:783] f, output logic [0:1411] leaf);
	assign leaf[0] = !f[358] && !f[357] && !f[359] && !f[384]; // c0t0i0
	assign leaf[1] = !f[358] && !f[357] && !f[359] && f[384]; // c0t0i0
	assign leaf[2] = !f[358] && !f[357] && f[359] && !f[462]; // c0t0i0
	assign leaf[3] = !f[358] && !f[357] && f[359] && f[462]; // c0t0i0
	assign leaf[4] = !f[358] && f[357] && !f[435] && !f[512]; // c0t0i0
	assign leaf[5] = !f[358] && f[357] && !f[435] && f[512]; // c0t0i0
	assign leaf[6] = !f[358] && f[357] && f[435] && !f[322]; // c0t0i0
	assign leaf[7] = !f[358] && f[357] && f[435] && f[322]; // c0t0i0
	assign leaf[8] = f[358] && !f[435] && !f[596] && !f[213]; // c0t0i0
	assign leaf[9] = f[358] && !f[435] && !f[596] && f[213]; // c0t0i0
	assign leaf[10] = f[358] && !f[435] && f[596] && !f[461]; // c0t0i0
	assign leaf[11] = f[358] && !f[435] && f[596] && f[461]; // c0t0i0
	assign leaf[12] = f[358] && f[435] && !f[295] && !f[245]; // c0t0i0
	assign leaf[13] = f[358] && f[435] && !f[295] && f[245]; // c0t0i0
	assign leaf[14] = f[358] && f[435] && f[295] && !f[538]; // c0t0i0
	assign leaf[15] = f[358] && f[435] && f[295] && f[538]; // c0t0i0
	assign leaf[16] = !f[407] && !f[463] && !f[351] && !f[627]; // c0t10i1
	assign leaf[17] = !f[407] && !f[463] && !f[351] && f[627]; // c0t10i1
	assign leaf[18] = !f[407] && !f[463] && f[351] && !f[455]; // c0t10i1
	assign leaf[19] = !f[407] && !f[463] && f[351] && f[455]; // c0t10i1
	assign leaf[20] = !f[407] && f[463] && !f[321] && !f[415]; // c0t10i1
	assign leaf[21] = !f[407] && f[463] && !f[321] && f[415]; // c0t10i1
	assign leaf[22] = !f[407] && f[463] && f[321] && !f[511]; // c0t10i1
	assign leaf[23] = !f[407] && f[463] && f[321] && f[511]; // c0t10i1
	assign leaf[24] = f[407] && !f[359] && !f[512]; // c0t10i1
	assign leaf[25] = f[407] && !f[359] && f[512] && !f[322]; // c0t10i1
	assign leaf[26] = f[407] && !f[359] && f[512] && f[322]; // c0t10i1
	assign leaf[27] = f[407] && f[359] && !f[509] && !f[188]; // c0t10i1
	assign leaf[28] = f[407] && f[359] && !f[509] && f[188]; // c0t10i1
	assign leaf[29] = f[407] && f[359] && f[509] && !f[296]; // c0t10i1
	assign leaf[30] = f[407] && f[359] && f[509] && f[296]; // c0t10i1
	assign leaf[31] = !f[407] && !f[490] && !f[352] && !f[184]; // c0t20i2
	assign leaf[32] = !f[407] && !f[490] && !f[352] && f[184]; // c0t20i2
	assign leaf[33] = !f[407] && !f[490] && f[352] && !f[456]; // c0t20i2
	assign leaf[34] = !f[407] && !f[490] && f[352] && f[456]; // c0t20i2
	assign leaf[35] = !f[407] && f[490] && !f[359] && !f[347]; // c0t20i2
	assign leaf[36] = !f[407] && f[490] && !f[359] && f[347]; // c0t20i2
	assign leaf[37] = !f[407] && f[490] && f[359] && !f[453]; // c0t20i2
	assign leaf[38] = !f[407] && f[490] && f[359] && f[453]; // c0t20i2
	assign leaf[39] = f[407] && !f[359] && !f[512]; // c0t20i2
	assign leaf[40] = f[407] && !f[359] && f[512] && !f[294]; // c0t20i2
	assign leaf[41] = f[407] && !f[359] && f[512] && f[294]; // c0t20i2
	assign leaf[42] = f[407] && f[359] && !f[322] && !f[187]; // c0t20i2
	assign leaf[43] = f[407] && f[359] && !f[322] && f[187]; // c0t20i2
	assign leaf[44] = f[407] && f[359] && f[322] && !f[432]; // c0t20i2
	assign leaf[45] = f[407] && f[359] && f[322] && f[432]; // c0t20i2
	assign leaf[46] = !f[434] && !f[380] && !f[489] && !f[484]; // c0t30i3
	assign leaf[47] = !f[434] && !f[380] && !f[489] && f[484]; // c0t30i3
	assign leaf[48] = !f[434] && !f[380] && f[489] && !f[386]; // c0t30i3
	assign leaf[49] = !f[434] && !f[380] && f[489] && f[386]; // c0t30i3
	assign leaf[50] = !f[434] && f[380] && !f[513] && !f[331]; // c0t30i3
	assign leaf[51] = !f[434] && f[380] && !f[513] && f[331]; // c0t30i3
	assign leaf[52] = !f[434] && f[380] && f[513] && !f[267]; // c0t30i3
	assign leaf[53] = !f[434] && f[380] && f[513] && f[267]; // c0t30i3
	assign leaf[54] = f[434] && !f[386] && !f[387]; // c0t30i3
	assign leaf[55] = f[434] && !f[386] && f[387] && !f[209]; // c0t30i3
	assign leaf[56] = f[434] && !f[386] && f[387] && f[209]; // c0t30i3
	assign leaf[57] = f[434] && f[386] && !f[625] && !f[219]; // c0t30i3
	assign leaf[58] = f[434] && f[386] && !f[625] && f[219]; // c0t30i3
	assign leaf[59] = f[434] && f[386] && f[625] && !f[468]; // c0t30i3
	assign leaf[60] = f[434] && f[386] && f[625] && f[468]; // c0t30i3
	assign leaf[61] = !f[407] && !f[511] && !f[513] && !f[481]; // c0t40i4
	assign leaf[62] = !f[407] && !f[511] && !f[513] && f[481]; // c0t40i4
	assign leaf[63] = !f[407] && !f[511] && f[513] && !f[490]; // c0t40i4
	assign leaf[64] = !f[407] && !f[511] && f[513] && f[490]; // c0t40i4
	assign leaf[65] = !f[407] && f[511] && !f[488] && !f[379]; // c0t40i4
	assign leaf[66] = !f[407] && f[511] && !f[488] && f[379]; // c0t40i4
	assign leaf[67] = !f[407] && f[511] && f[488] && !f[400]; // c0t40i4
	assign leaf[68] = !f[407] && f[511] && f[488] && f[400]; // c0t40i4
	assign leaf[69] = f[407] && !f[359] && !f[512] && !f[396]; // c0t40i4
	assign leaf[70] = f[407] && !f[359] && !f[512] && f[396]; // c0t40i4
	assign leaf[71] = f[407] && !f[359] && f[512] && !f[655]; // c0t40i4
	assign leaf[72] = f[407] && !f[359] && f[512] && f[655]; // c0t40i4
	assign leaf[73] = f[407] && f[359] && !f[245] && !f[453]; // c0t40i4
	assign leaf[74] = f[407] && f[359] && !f[245] && f[453]; // c0t40i4
	assign leaf[75] = f[407] && f[359] && f[245] && !f[468]; // c0t40i4
	assign leaf[76] = f[407] && f[359] && f[245] && f[468]; // c0t40i4
	assign leaf[77] = !f[435] && !f[379] && !f[598] && !f[539]; // c0t50i5
	assign leaf[78] = !f[435] && !f[379] && !f[598] && f[539]; // c0t50i5
	assign leaf[79] = !f[435] && !f[379] && f[598] && !f[489]; // c0t50i5
	assign leaf[80] = !f[435] && !f[379] && f[598] && f[489]; // c0t50i5
	assign leaf[81] = !f[435] && f[379] && !f[331] && !f[329]; // c0t50i5
	assign leaf[82] = !f[435] && f[379] && !f[331] && f[329]; // c0t50i5
	assign leaf[83] = !f[435] && f[379] && f[331] && !f[265]; // c0t50i5
	assign leaf[84] = !f[435] && f[379] && f[331] && f[265]; // c0t50i5
	assign leaf[85] = f[435] && !f[386] && !f[540] && !f[539]; // c0t50i5
	assign leaf[86] = f[435] && !f[386] && !f[540] && f[539]; // c0t50i5
	assign leaf[87] = f[435] && !f[386] && f[540] && !f[434]; // c0t50i5
	assign leaf[88] = f[435] && !f[386] && f[540] && f[434]; // c0t50i5
	assign leaf[89] = f[435] && f[386] && !f[322] && !f[625]; // c0t50i5
	assign leaf[90] = f[435] && f[386] && !f[322] && f[625]; // c0t50i5
	assign leaf[91] = f[435] && f[386] && f[322] && !f[433]; // c0t50i5
	assign leaf[92] = f[435] && f[386] && f[322] && f[433]; // c0t50i5
	assign leaf[93] = !f[434] && !f[455] && !f[457] && !f[425]; // c0t60i6
	assign leaf[94] = !f[434] && !f[455] && !f[457] && f[425]; // c0t60i6
	assign leaf[95] = !f[434] && !f[455] && f[457] && !f[628]; // c0t60i6
	assign leaf[96] = !f[434] && !f[455] && f[457] && f[628]; // c0t60i6
	assign leaf[97] = !f[434] && f[455] && !f[626] && !f[410]; // c0t60i6
	assign leaf[98] = !f[434] && f[455] && !f[626] && f[410]; // c0t60i6
	assign leaf[99] = !f[434] && f[455] && f[626] && !f[378]; // c0t60i6
	assign leaf[100] = !f[434] && f[455] && f[626] && f[378]; // c0t60i6
	assign leaf[101] = f[434] && !f[385] && !f[359]; // c0t60i6
	assign leaf[102] = f[434] && !f[385] && f[359] && !f[185]; // c0t60i6
	assign leaf[103] = f[434] && !f[385] && f[359] && f[185]; // c0t60i6
	assign leaf[104] = f[434] && f[385] && !f[409] && !f[655]; // c0t60i6
	assign leaf[105] = f[434] && f[385] && !f[409] && f[655]; // c0t60i6
	assign leaf[106] = f[434] && f[385] && f[409] && !f[274]; // c0t60i6
	assign leaf[107] = f[434] && f[385] && f[409] && f[274]; // c0t60i6
	assign leaf[108] = !f[408] && !f[461] && !f[352] && !f[214]; // c0t70i7
	assign leaf[109] = !f[408] && !f[461] && !f[352] && f[214]; // c0t70i7
	assign leaf[110] = !f[408] && !f[461] && f[352] && !f[265]; // c0t70i7
	assign leaf[111] = !f[408] && !f[461] && f[352] && f[265]; // c0t70i7
	assign leaf[112] = !f[408] && f[461] && !f[386] && !f[657]; // c0t70i7
	assign leaf[113] = !f[408] && f[461] && !f[386] && f[657]; // c0t70i7
	assign leaf[114] = !f[408] && f[461] && f[386] && !f[293]; // c0t70i7
	assign leaf[115] = !f[408] && f[461] && f[386] && f[293]; // c0t70i7
	assign leaf[116] = f[408] && !f[484] && !f[514] && !f[481]; // c0t70i7
	assign leaf[117] = f[408] && !f[484] && !f[514] && f[481]; // c0t70i7
	assign leaf[118] = f[408] && !f[484] && f[514] && !f[434]; // c0t70i7
	assign leaf[119] = f[408] && !f[484] && f[514] && f[434]; // c0t70i7
	assign leaf[120] = f[408] && f[484] && !f[626] && !f[331]; // c0t70i7
	assign leaf[121] = f[408] && f[484] && !f[626] && f[331]; // c0t70i7
	assign leaf[122] = f[408] && f[484] && f[626] && !f[433]; // c0t70i7
	assign leaf[123] = f[408] && f[484] && f[626] && f[433]; // c0t70i7
	assign leaf[124] = !f[408] && !f[427] && !f[429] && !f[425]; // c0t80i8
	assign leaf[125] = !f[408] && !f[427] && !f[429] && f[425]; // c0t80i8
	assign leaf[126] = !f[408] && !f[427] && f[429] && !f[485]; // c0t80i8
	assign leaf[127] = !f[408] && !f[427] && f[429] && f[485]; // c0t80i8
	assign leaf[128] = !f[408] && f[427] && !f[460] && !f[716]; // c0t80i8
	assign leaf[129] = !f[408] && f[427] && !f[460] && f[716]; // c0t80i8
	assign leaf[130] = !f[408] && f[427] && f[460] && !f[292]; // c0t80i8
	assign leaf[131] = !f[408] && f[427] && f[460] && f[292]; // c0t80i8
	assign leaf[132] = f[408] && !f[293] && !f[455]; // c0t80i8
	assign leaf[133] = f[408] && !f[293] && f[455] && !f[656]; // c0t80i8
	assign leaf[134] = f[408] && !f[293] && f[455] && f[656]; // c0t80i8
	assign leaf[135] = f[408] && f[293] && !f[406] && !f[404]; // c0t80i8
	assign leaf[136] = f[408] && f[293] && !f[406] && f[404]; // c0t80i8
	assign leaf[137] = f[408] && f[293] && f[406] && !f[414]; // c0t80i8
	assign leaf[138] = f[408] && f[293] && f[406] && f[414]; // c0t80i8
	assign leaf[139] = !f[462] && !f[378] && !f[402] && !f[410]; // c0t90i9
	assign leaf[140] = !f[462] && !f[378] && !f[402] && f[410]; // c0t90i9
	assign leaf[141] = !f[462] && !f[378] && f[402] && !f[599]; // c0t90i9
	assign leaf[142] = !f[462] && !f[378] && f[402] && f[599]; // c0t90i9
	assign leaf[143] = !f[462] && f[378] && !f[273] && !f[274]; // c0t90i9
	assign leaf[144] = !f[462] && f[378] && !f[273] && f[274]; // c0t90i9
	assign leaf[145] = !f[462] && f[378] && f[273] && !f[266]; // c0t90i9
	assign leaf[146] = !f[462] && f[378] && f[273] && f[266]; // c0t90i9
	assign leaf[147] = f[462] && !f[386] && !f[568] && !f[508]; // c0t90i9
	assign leaf[148] = f[462] && !f[386] && !f[568] && f[508]; // c0t90i9
	assign leaf[149] = f[462] && !f[386] && f[568] && !f[461]; // c0t90i9
	assign leaf[150] = f[462] && !f[386] && f[568] && f[461]; // c0t90i9
	assign leaf[151] = f[462] && f[386] && !f[297] && !f[273]; // c0t90i9
	assign leaf[152] = f[462] && f[386] && !f[297] && f[273]; // c0t90i9
	assign leaf[153] = f[462] && f[386] && f[297] && !f[155]; // c0t90i9
	assign leaf[154] = f[462] && f[386] && f[297] && f[155]; // c0t90i9
	assign leaf[155] = !f[434] && !f[455] && !f[458] && !f[425]; // c0t100i10
	assign leaf[156] = !f[434] && !f[455] && !f[458] && f[425]; // c0t100i10
	assign leaf[157] = !f[434] && !f[455] && f[458] && !f[355]; // c0t100i10
	assign leaf[158] = !f[434] && !f[455] && f[458] && f[355]; // c0t100i10
	assign leaf[159] = !f[434] && f[455] && !f[539] && !f[437]; // c0t100i10
	assign leaf[160] = !f[434] && f[455] && !f[539] && f[437]; // c0t100i10
	assign leaf[161] = !f[434] && f[455] && f[539] && !f[98]; // c0t100i10
	assign leaf[162] = !f[434] && f[455] && f[539] && f[98]; // c0t100i10
	assign leaf[163] = f[434] && !f[385] && !f[360] && !f[383]; // c0t100i10
	assign leaf[164] = f[434] && !f[385] && !f[360] && f[383]; // c0t100i10
	assign leaf[165] = f[434] && !f[385] && f[360]; // c0t100i10
	assign leaf[166] = f[434] && f[385] && !f[468] && !f[536]; // c0t100i10
	assign leaf[167] = f[434] && f[385] && !f[468] && f[536]; // c0t100i10
	assign leaf[168] = f[434] && f[385] && f[468] && !f[213]; // c0t100i10
	assign leaf[169] = f[434] && f[385] && f[468] && f[213]; // c0t100i10
	assign leaf[170] = !f[379] && !f[491] && !f[323] && !f[436]; // c0t110i11
	assign leaf[171] = !f[379] && !f[491] && !f[323] && f[436]; // c0t110i11
	assign leaf[172] = !f[379] && !f[491] && f[323] && !f[239]; // c0t110i11
	assign leaf[173] = !f[379] && !f[491] && f[323] && f[239]; // c0t110i11
	assign leaf[174] = !f[379] && f[491] && !f[348] && !f[387]; // c0t110i11
	assign leaf[175] = !f[379] && f[491] && !f[348] && f[387]; // c0t110i11
	assign leaf[176] = !f[379] && f[491] && f[348] && !f[625]; // c0t110i11
	assign leaf[177] = !f[379] && f[491] && f[348] && f[625]; // c0t110i11
	assign leaf[178] = f[379] && !f[329] && !f[331] && !f[513]; // c0t110i11
	assign leaf[179] = f[379] && !f[329] && !f[331] && f[513]; // c0t110i11
	assign leaf[180] = f[379] && !f[329] && f[331] && !f[346]; // c0t110i11
	assign leaf[181] = f[379] && !f[329] && f[331] && f[346]; // c0t110i11
	assign leaf[182] = f[379] && f[329] && !f[215] && !f[443]; // c0t110i11
	assign leaf[183] = f[379] && f[329] && !f[215] && f[443]; // c0t110i11
	assign leaf[184] = f[379] && f[329] && f[215] && !f[382]; // c0t110i11
	assign leaf[185] = f[379] && f[329] && f[215] && f[382]; // c0t110i11
	assign leaf[186] = !f[387] && !f[429] && !f[427] && !f[430]; // c0t120i12
	assign leaf[187] = !f[387] && !f[429] && !f[427] && f[430]; // c0t120i12
	assign leaf[188] = !f[387] && !f[429] && f[427] && !f[625]; // c0t120i12
	assign leaf[189] = !f[387] && !f[429] && f[427] && f[625]; // c0t120i12
	assign leaf[190] = !f[387] && f[429] && !f[627] && !f[624]; // c0t120i12
	assign leaf[191] = !f[387] && f[429] && !f[627] && f[624]; // c0t120i12
	assign leaf[192] = !f[387] && f[429] && f[627] && !f[513]; // c0t120i12
	assign leaf[193] = !f[387] && f[429] && f[627] && f[513]; // c0t120i12
	assign leaf[194] = f[387] && !f[426] && !f[302] && !f[304]; // c0t120i12
	assign leaf[195] = f[387] && !f[426] && !f[302] && f[304]; // c0t120i12
	assign leaf[196] = f[387] && !f[426] && f[302] && !f[539]; // c0t120i12
	assign leaf[197] = f[387] && !f[426] && f[302] && f[539]; // c0t120i12
	assign leaf[198] = f[387] && f[426] && !f[437] && !f[433]; // c0t120i12
	assign leaf[199] = f[387] && f[426] && !f[437] && f[433]; // c0t120i12
	assign leaf[200] = f[387] && f[426] && f[437] && !f[301]; // c0t120i12
	assign leaf[201] = f[387] && f[426] && f[437] && f[301]; // c0t120i12
	assign leaf[202] = !f[434] && !f[242] && !f[387] && !f[240]; // c0t130i13
	assign leaf[203] = !f[434] && !f[242] && !f[387] && f[240]; // c0t130i13
	assign leaf[204] = !f[434] && !f[242] && f[387] && !f[350]; // c0t130i13
	assign leaf[205] = !f[434] && !f[242] && f[387] && f[350]; // c0t130i13
	assign leaf[206] = !f[434] && f[242] && !f[570] && !f[624]; // c0t130i13
	assign leaf[207] = !f[434] && f[242] && !f[570] && f[624]; // c0t130i13
	assign leaf[208] = !f[434] && f[242] && f[570] && !f[401]; // c0t130i13
	assign leaf[209] = !f[434] && f[242] && f[570] && f[401]; // c0t130i13
	assign leaf[210] = f[434] && !f[540] && !f[537]; // c0t130i13
	assign leaf[211] = f[434] && !f[540] && f[537] && !f[323]; // c0t130i13
	assign leaf[212] = f[434] && !f[540] && f[537] && f[323]; // c0t130i13
	assign leaf[213] = f[434] && f[540] && !f[344] && !f[374]; // c0t130i13
	assign leaf[214] = f[434] && f[540] && !f[344] && f[374]; // c0t130i13
	assign leaf[215] = f[434] && f[540] && f[344] && !f[656]; // c0t130i13
	assign leaf[216] = f[434] && f[540] && f[344] && f[656]; // c0t130i13
	assign leaf[217] = !f[406] && !f[490] && !f[323] && !f[629]; // c0t140i14
	assign leaf[218] = !f[406] && !f[490] && !f[323] && f[629]; // c0t140i14
	assign leaf[219] = !f[406] && !f[490] && f[323] && !f[239]; // c0t140i14
	assign leaf[220] = !f[406] && !f[490] && f[323] && f[239]; // c0t140i14
	assign leaf[221] = !f[406] && f[490] && !f[294] && !f[415]; // c0t140i14
	assign leaf[222] = !f[406] && f[490] && !f[294] && f[415]; // c0t140i14
	assign leaf[223] = !f[406] && f[490] && f[294] && !f[570]; // c0t140i14
	assign leaf[224] = !f[406] && f[490] && f[294] && f[570]; // c0t140i14
	assign leaf[225] = f[406] && !f[329] && !f[332] && !f[328]; // c0t140i14
	assign leaf[226] = f[406] && !f[329] && !f[332] && f[328]; // c0t140i14
	assign leaf[227] = f[406] && !f[329] && f[332] && !f[656]; // c0t140i14
	assign leaf[228] = f[406] && !f[329] && f[332] && f[656]; // c0t140i14
	assign leaf[229] = f[406] && f[329] && !f[295] && !f[404]; // c0t140i14
	assign leaf[230] = f[406] && f[329] && !f[295] && f[404]; // c0t140i14
	assign leaf[231] = f[406] && f[329] && f[295] && !f[412]; // c0t140i14
	assign leaf[232] = f[406] && f[329] && f[295] && f[412]; // c0t140i14
	assign leaf[233] = !f[379] && !f[491] && !f[322] && !f[435]; // c0t150i15
	assign leaf[234] = !f[379] && !f[491] && !f[322] && f[435]; // c0t150i15
	assign leaf[235] = !f[379] && !f[491] && f[322] && !f[273]; // c0t150i15
	assign leaf[236] = !f[379] && !f[491] && f[322] && f[273]; // c0t150i15
	assign leaf[237] = !f[379] && f[491] && !f[348] && !f[415]; // c0t150i15
	assign leaf[238] = !f[379] && f[491] && !f[348] && f[415]; // c0t150i15
	assign leaf[239] = !f[379] && f[491] && f[348] && !f[598]; // c0t150i15
	assign leaf[240] = !f[379] && f[491] && f[348] && f[598]; // c0t150i15
	assign leaf[241] = f[379] && !f[329] && !f[331] && !f[486]; // c0t150i15
	assign leaf[242] = f[379] && !f[329] && !f[331] && f[486]; // c0t150i15
	assign leaf[243] = f[379] && !f[329] && f[331] && !f[604]; // c0t150i15
	assign leaf[244] = f[379] && !f[329] && f[331] && f[604]; // c0t150i15
	assign leaf[245] = f[379] && f[329] && !f[268] && !f[431]; // c0t150i15
	assign leaf[246] = f[379] && f[329] && !f[268] && f[431]; // c0t150i15
	assign leaf[247] = f[379] && f[329] && f[268] && !f[540]; // c0t150i15
	assign leaf[248] = f[379] && f[329] && f[268] && f[540]; // c0t150i15
	assign leaf[249] = !f[482] && !f[485] && !f[486] && !f[480]; // c0t160i16
	assign leaf[250] = !f[482] && !f[485] && !f[486] && f[480]; // c0t160i16
	assign leaf[251] = !f[482] && !f[485] && f[486] && !f[154]; // c0t160i16
	assign leaf[252] = !f[482] && !f[485] && f[486] && f[154]; // c0t160i16
	assign leaf[253] = !f[482] && f[485] && !f[656] && !f[600]; // c0t160i16
	assign leaf[254] = !f[482] && f[485] && !f[656] && f[600]; // c0t160i16
	assign leaf[255] = !f[482] && f[485] && f[656] && !f[541]; // c0t160i16
	assign leaf[256] = !f[482] && f[485] && f[656] && f[541]; // c0t160i16
	assign leaf[257] = f[482] && !f[399] && !f[516] && !f[462]; // c0t160i16
	assign leaf[258] = f[482] && !f[399] && !f[516] && f[462]; // c0t160i16
	assign leaf[259] = f[482] && !f[399] && f[516] && !f[219]; // c0t160i16
	assign leaf[260] = f[482] && !f[399] && f[516] && f[219]; // c0t160i16
	assign leaf[261] = f[482] && f[399] && !f[409] && !f[691]; // c0t160i16
	assign leaf[262] = f[482] && f[399] && !f[409] && f[691]; // c0t160i16
	assign leaf[263] = f[482] && f[399] && f[409] && !f[320]; // c0t160i16
	assign leaf[264] = f[482] && f[399] && f[409] && f[320]; // c0t160i16
	assign leaf[265] = !f[406] && !f[387] && !f[402] && !f[400]; // c0t170i17
	assign leaf[266] = !f[406] && !f[387] && !f[402] && f[400]; // c0t170i17
	assign leaf[267] = !f[406] && !f[387] && f[402] && !f[299]; // c0t170i17
	assign leaf[268] = !f[406] && !f[387] && f[402] && f[299]; // c0t170i17
	assign leaf[269] = !f[406] && f[387] && !f[510] && !f[398]; // c0t170i17
	assign leaf[270] = !f[406] && f[387] && !f[510] && f[398]; // c0t170i17
	assign leaf[271] = !f[406] && f[387] && f[510] && !f[437]; // c0t170i17
	assign leaf[272] = !f[406] && f[387] && f[510] && f[437]; // c0t170i17
	assign leaf[273] = f[406] && !f[244] && !f[405] && !f[356]; // c0t170i17
	assign leaf[274] = f[406] && !f[244] && !f[405] && f[356]; // c0t170i17
	assign leaf[275] = f[406] && !f[244] && f[405] && !f[621]; // c0t170i17
	assign leaf[276] = f[406] && !f[244] && f[405] && f[621]; // c0t170i17
	assign leaf[277] = f[406] && f[244] && !f[540] && !f[508]; // c0t170i17
	assign leaf[278] = f[406] && f[244] && !f[540] && f[508]; // c0t170i17
	assign leaf[279] = f[406] && f[244] && f[540] && !f[357]; // c0t170i17
	assign leaf[280] = f[406] && f[244] && f[540] && f[357]; // c0t170i17
	assign leaf[281] = !f[379] && !f[518] && !f[323] && !f[462]; // c0t180i18
	assign leaf[282] = !f[379] && !f[518] && !f[323] && f[462]; // c0t180i18
	assign leaf[283] = !f[379] && !f[518] && f[323] && !f[238]; // c0t180i18
	assign leaf[284] = !f[379] && !f[518] && f[323] && f[238]; // c0t180i18
	assign leaf[285] = !f[379] && f[518] && !f[321] && !f[387]; // c0t180i18
	assign leaf[286] = !f[379] && f[518] && !f[321] && f[387]; // c0t180i18
	assign leaf[287] = !f[379] && f[518] && f[321] && !f[427]; // c0t180i18
	assign leaf[288] = !f[379] && f[518] && f[321] && f[427]; // c0t180i18
	assign leaf[289] = f[379] && !f[569] && !f[293] && !f[541]; // c0t180i18
	assign leaf[290] = f[379] && !f[569] && !f[293] && f[541]; // c0t180i18
	assign leaf[291] = f[379] && !f[569] && f[293] && !f[576]; // c0t180i18
	assign leaf[292] = f[379] && !f[569] && f[293] && f[576]; // c0t180i18
	assign leaf[293] = f[379] && f[569] && !f[377] && !f[656]; // c0t180i18
	assign leaf[294] = f[379] && f[569] && !f[377] && f[656]; // c0t180i18
	assign leaf[295] = f[379] && f[569] && f[377] && !f[380]; // c0t180i18
	assign leaf[296] = f[379] && f[569] && f[377] && f[380]; // c0t180i18
	assign leaf[297] = !f[570] && !f[624] && !f[543] && !f[623]; // c0t190i19
	assign leaf[298] = !f[570] && !f[624] && !f[543] && f[623]; // c0t190i19
	assign leaf[299] = !f[570] && !f[624] && f[543] && !f[491]; // c0t190i19
	assign leaf[300] = !f[570] && !f[624] && f[543] && f[491]; // c0t190i19
	assign leaf[301] = !f[570] && f[624] && !f[152] && !f[487]; // c0t190i19
	assign leaf[302] = !f[570] && f[624] && !f[152] && f[487]; // c0t190i19
	assign leaf[303] = !f[570] && f[624] && f[152] && !f[397]; // c0t190i19
	assign leaf[304] = !f[570] && f[624] && f[152] && f[397]; // c0t190i19
	assign leaf[305] = f[570] && !f[656] && !f[371] && !f[401]; // c0t190i19
	assign leaf[306] = f[570] && !f[656] && !f[371] && f[401]; // c0t190i19
	assign leaf[307] = f[570] && !f[656] && f[371] && !f[265]; // c0t190i19
	assign leaf[308] = f[570] && !f[656] && f[371] && f[265]; // c0t190i19
	assign leaf[309] = f[570] && f[656] && !f[486] && !f[456]; // c0t190i19
	assign leaf[310] = f[570] && f[656] && !f[486] && f[456]; // c0t190i19
	assign leaf[311] = f[570] && f[656] && f[486] && !f[608]; // c0t190i19
	assign leaf[312] = f[570] && f[656] && f[486] && f[608]; // c0t190i19
	assign leaf[313] = !f[415] && !f[401] && !f[403] && !f[399]; // c0t200i20
	assign leaf[314] = !f[415] && !f[401] && !f[403] && f[399]; // c0t200i20
	assign leaf[315] = !f[415] && !f[401] && f[403] && !f[514]; // c0t200i20
	assign leaf[316] = !f[415] && !f[401] && f[403] && f[514]; // c0t200i20
	assign leaf[317] = !f[415] && f[401] && !f[484] && !f[542]; // c0t200i20
	assign leaf[318] = !f[415] && f[401] && !f[484] && f[542]; // c0t200i20
	assign leaf[319] = !f[415] && f[401] && f[484] && !f[654]; // c0t200i20
	assign leaf[320] = !f[415] && f[401] && f[484] && f[654]; // c0t200i20
	assign leaf[321] = f[415] && !f[425] && !f[275] && !f[302]; // c0t200i20
	assign leaf[322] = f[415] && !f[425] && !f[275] && f[302]; // c0t200i20
	assign leaf[323] = f[415] && !f[425] && f[275] && !f[319]; // c0t200i20
	assign leaf[324] = f[415] && !f[425] && f[275] && f[319]; // c0t200i20
	assign leaf[325] = f[415] && f[425] && !f[404] && !f[148]; // c0t200i20
	assign leaf[326] = f[415] && f[425] && !f[404] && f[148]; // c0t200i20
	assign leaf[327] = f[415] && f[425] && f[404] && !f[346]; // c0t200i20
	assign leaf[328] = f[415] && f[425] && f[404] && f[346]; // c0t200i20
	assign leaf[329] = !f[240] && !f[350] && !f[518] && !f[214]; // c0t210i21
	assign leaf[330] = !f[240] && !f[350] && !f[518] && f[214]; // c0t210i21
	assign leaf[331] = !f[240] && !f[350] && f[518] && !f[442]; // c0t210i21
	assign leaf[332] = !f[240] && !f[350] && f[518] && f[442]; // c0t210i21
	assign leaf[333] = !f[240] && f[350] && !f[215] && !f[190]; // c0t210i21
	assign leaf[334] = !f[240] && f[350] && !f[215] && f[190]; // c0t210i21
	assign leaf[335] = !f[240] && f[350] && f[215] && !f[264]; // c0t210i21
	assign leaf[336] = !f[240] && f[350] && f[215] && f[264]; // c0t210i21
	assign leaf[337] = f[240] && !f[462] && !f[690] && !f[712]; // c0t210i21
	assign leaf[338] = f[240] && !f[462] && !f[690] && f[712]; // c0t210i21
	assign leaf[339] = f[240] && !f[462] && f[690] && !f[498]; // c0t210i21
	assign leaf[340] = f[240] && !f[462] && f[690] && f[498]; // c0t210i21
	assign leaf[341] = f[240] && f[462] && !f[512] && !f[480]; // c0t210i21
	assign leaf[342] = f[240] && f[462] && !f[512] && f[480]; // c0t210i21
	assign leaf[343] = f[240] && f[462] && f[512] && !f[401]; // c0t210i21
	assign leaf[344] = f[240] && f[462] && f[512] && f[401]; // c0t210i21
	assign leaf[345] = !f[453] && !f[429] && !f[431] && !f[427]; // c0t220i22
	assign leaf[346] = !f[453] && !f[429] && !f[431] && f[427]; // c0t220i22
	assign leaf[347] = !f[453] && !f[429] && f[431] && !f[241]; // c0t220i22
	assign leaf[348] = !f[453] && !f[429] && f[431] && f[241]; // c0t220i22
	assign leaf[349] = !f[453] && f[429] && !f[513] && !f[511]; // c0t220i22
	assign leaf[350] = !f[453] && f[429] && !f[513] && f[511]; // c0t220i22
	assign leaf[351] = !f[453] && f[429] && f[513] && !f[328]; // c0t220i22
	assign leaf[352] = !f[453] && f[429] && f[513] && f[328]; // c0t220i22
	assign leaf[353] = f[453] && !f[458] && !f[623] && !f[410]; // c0t220i22
	assign leaf[354] = f[453] && !f[458] && !f[623] && f[410]; // c0t220i22
	assign leaf[355] = f[453] && !f[458] && f[623] && !f[404]; // c0t220i22
	assign leaf[356] = f[453] && !f[458] && f[623] && f[404]; // c0t220i22
	assign leaf[357] = f[453] && f[458] && !f[346] && !f[470]; // c0t220i22
	assign leaf[358] = f[453] && f[458] && !f[346] && f[470]; // c0t220i22
	assign leaf[359] = f[453] && f[458] && f[346] && !f[544]; // c0t220i22
	assign leaf[360] = f[453] && f[458] && f[346] && f[544]; // c0t220i22
	assign leaf[361] = !f[663] && !f[434] && !f[241] && !f[215]; // c0t230i23
	assign leaf[362] = !f[663] && !f[434] && !f[241] && f[215]; // c0t230i23
	assign leaf[363] = !f[663] && !f[434] && f[241] && !f[713]; // c0t230i23
	assign leaf[364] = !f[663] && !f[434] && f[241] && f[713]; // c0t230i23
	assign leaf[365] = !f[663] && f[434] && !f[540] && !f[481]; // c0t230i23
	assign leaf[366] = !f[663] && f[434] && !f[540] && f[481]; // c0t230i23
	assign leaf[367] = !f[663] && f[434] && f[540] && !f[328]; // c0t230i23
	assign leaf[368] = !f[663] && f[434] && f[540] && f[328]; // c0t230i23
	assign leaf[369] = f[663] && !f[526] && !f[546] && !f[572]; // c0t230i23
	assign leaf[370] = f[663] && !f[526] && !f[546] && f[572]; // c0t230i23
	assign leaf[371] = f[663] && !f[526] && f[546] && !f[464]; // c0t230i23
	assign leaf[372] = f[663] && !f[526] && f[546] && f[464]; // c0t230i23
	assign leaf[373] = f[663] && f[526] && !f[347] && !f[402]; // c0t230i23
	assign leaf[374] = f[663] && f[526] && !f[347] && f[402]; // c0t230i23
	assign leaf[375] = f[663] && f[526] && f[347] && !f[551]; // c0t230i23
	assign leaf[376] = f[663] && f[526] && f[347] && f[551]; // c0t230i23
	assign leaf[377] = !f[663] && !f[406] && !f[688] && !f[398]; // c0t240i24
	assign leaf[378] = !f[663] && !f[406] && !f[688] && f[398]; // c0t240i24
	assign leaf[379] = !f[663] && !f[406] && f[688] && !f[656]; // c0t240i24
	assign leaf[380] = !f[663] && !f[406] && f[688] && f[656]; // c0t240i24
	assign leaf[381] = !f[663] && f[406] && !f[380] && !f[347]; // c0t240i24
	assign leaf[382] = !f[663] && f[406] && !f[380] && f[347]; // c0t240i24
	assign leaf[383] = !f[663] && f[406] && f[380] && !f[571]; // c0t240i24
	assign leaf[384] = !f[663] && f[406] && f[380] && f[571]; // c0t240i24
	assign leaf[385] = f[663] && !f[526] && !f[687] && !f[638]; // c0t240i24
	assign leaf[386] = f[663] && !f[526] && !f[687] && f[638]; // c0t240i24
	assign leaf[387] = f[663] && !f[526] && f[687] && !f[204]; // c0t240i24
	assign leaf[388] = f[663] && !f[526] && f[687] && f[204]; // c0t240i24
	assign leaf[389] = f[663] && f[526] && !f[347] && !f[402]; // c0t240i24
	assign leaf[390] = f[663] && f[526] && !f[347] && f[402]; // c0t240i24
	assign leaf[391] = f[663] && f[526] && f[347] && !f[572]; // c0t240i24
	assign leaf[392] = f[663] && f[526] && f[347] && f[572]; // c0t240i24
	assign leaf[393] = !f[434] && !f[177] && !f[517] && !f[350]; // c0t250i25
	assign leaf[394] = !f[434] && !f[177] && !f[517] && f[350]; // c0t250i25
	assign leaf[395] = !f[434] && !f[177] && f[517] && !f[297]; // c0t250i25
	assign leaf[396] = !f[434] && !f[177] && f[517] && f[297]; // c0t250i25
	assign leaf[397] = !f[434] && f[177] && !f[397] && !f[596]; // c0t250i25
	assign leaf[398] = !f[434] && f[177] && !f[397] && f[596]; // c0t250i25
	assign leaf[399] = !f[434] && f[177] && f[397] && !f[633]; // c0t250i25
	assign leaf[400] = !f[434] && f[177] && f[397] && f[633]; // c0t250i25
	assign leaf[401] = f[434] && !f[569] && !f[161]; // c0t250i25
	assign leaf[402] = f[434] && !f[569] && f[161]; // c0t250i25
	assign leaf[403] = f[434] && f[569] && !f[428] && !f[601]; // c0t250i25
	assign leaf[404] = f[434] && f[569] && !f[428] && f[601]; // c0t250i25
	assign leaf[405] = f[434] && f[569] && f[428] && !f[431]; // c0t250i25
	assign leaf[406] = f[434] && f[569] && f[428] && f[431]; // c0t250i25
	assign leaf[407] = !f[542] && !f[510] && !f[512] && !f[471]; // c0t260i26
	assign leaf[408] = !f[542] && !f[510] && !f[512] && f[471]; // c0t260i26
	assign leaf[409] = !f[542] && !f[510] && f[512] && !f[654]; // c0t260i26
	assign leaf[410] = !f[542] && !f[510] && f[512] && f[654]; // c0t260i26
	assign leaf[411] = !f[542] && f[510] && !f[246] && !f[404]; // c0t260i26
	assign leaf[412] = !f[542] && f[510] && !f[246] && f[404]; // c0t260i26
	assign leaf[413] = !f[542] && f[510] && f[246] && !f[487]; // c0t260i26
	assign leaf[414] = !f[542] && f[510] && f[246] && f[487]; // c0t260i26
	assign leaf[415] = f[542] && !f[298] && !f[272] && !f[297]; // c0t260i26
	assign leaf[416] = f[542] && !f[298] && !f[272] && f[297]; // c0t260i26
	assign leaf[417] = f[542] && !f[298] && f[272] && !f[545]; // c0t260i26
	assign leaf[418] = f[542] && !f[298] && f[272] && f[545]; // c0t260i26
	assign leaf[419] = f[542] && f[298] && !f[430] && !f[415]; // c0t260i26
	assign leaf[420] = f[542] && f[298] && !f[430] && f[415]; // c0t260i26
	assign leaf[421] = f[542] && f[298] && f[430] && !f[383]; // c0t260i26
	assign leaf[422] = f[542] && f[298] && f[430] && f[383]; // c0t260i26
	assign leaf[423] = !f[378] && !f[571] && !f[654] && !f[415]; // c0t270i27
	assign leaf[424] = !f[378] && !f[571] && !f[654] && f[415]; // c0t270i27
	assign leaf[425] = !f[378] && !f[571] && f[654] && !f[455]; // c0t270i27
	assign leaf[426] = !f[378] && !f[571] && f[654] && f[455]; // c0t270i27
	assign leaf[427] = !f[378] && f[571] && !f[681] && !f[159]; // c0t270i27
	assign leaf[428] = !f[378] && f[571] && !f[681] && f[159]; // c0t270i27
	assign leaf[429] = !f[378] && f[571] && f[681] && !f[511]; // c0t270i27
	assign leaf[430] = !f[378] && f[571] && f[681] && f[511]; // c0t270i27
	assign leaf[431] = f[378] && !f[294] && !f[376] && !f[496]; // c0t270i27
	assign leaf[432] = f[378] && !f[294] && !f[376] && f[496]; // c0t270i27
	assign leaf[433] = f[378] && !f[294] && f[376] && !f[353]; // c0t270i27
	assign leaf[434] = f[378] && !f[294] && f[376] && f[353]; // c0t270i27
	assign leaf[435] = f[378] && f[294] && !f[245] && !f[438]; // c0t270i27
	assign leaf[436] = f[378] && f[294] && !f[245] && f[438]; // c0t270i27
	assign leaf[437] = f[378] && f[294] && f[245] && !f[352]; // c0t270i27
	assign leaf[438] = f[378] && f[294] && f[245] && f[352]; // c0t270i27
	assign leaf[439] = !f[265] && !f[351] && !f[493] && !f[321]; // c0t280i28
	assign leaf[440] = !f[265] && !f[351] && !f[493] && f[321]; // c0t280i28
	assign leaf[441] = !f[265] && !f[351] && f[493] && !f[288]; // c0t280i28
	assign leaf[442] = !f[265] && !f[351] && f[493] && f[288]; // c0t280i28
	assign leaf[443] = !f[265] && f[351] && !f[216] && !f[347]; // c0t280i28
	assign leaf[444] = !f[265] && f[351] && !f[216] && f[347]; // c0t280i28
	assign leaf[445] = !f[265] && f[351] && f[216] && !f[353]; // c0t280i28
	assign leaf[446] = !f[265] && f[351] && f[216] && f[353]; // c0t280i28
	assign leaf[447] = f[265] && !f[416] && !f[347] && !f[469]; // c0t280i28
	assign leaf[448] = f[265] && !f[416] && !f[347] && f[469]; // c0t280i28
	assign leaf[449] = f[265] && !f[416] && f[347] && !f[635]; // c0t280i28
	assign leaf[450] = f[265] && !f[416] && f[347] && f[635]; // c0t280i28
	assign leaf[451] = f[265] && f[416] && !f[414]; // c0t280i28
	assign leaf[452] = f[265] && f[416] && f[414] && !f[398]; // c0t280i28
	assign leaf[453] = f[265] && f[416] && f[414] && f[398]; // c0t280i28
	assign leaf[454] = !f[663] && !f[453] && !f[486] && !f[456]; // c0t290i29
	assign leaf[455] = !f[663] && !f[453] && !f[486] && f[456]; // c0t290i29
	assign leaf[456] = !f[663] && !f[453] && f[486] && !f[489]; // c0t290i29
	assign leaf[457] = !f[663] && !f[453] && f[486] && f[489]; // c0t290i29
	assign leaf[458] = !f[663] && f[453] && !f[303] && !f[329]; // c0t290i29
	assign leaf[459] = !f[663] && f[453] && !f[303] && f[329]; // c0t290i29
	assign leaf[460] = !f[663] && f[453] && f[303] && !f[150]; // c0t290i29
	assign leaf[461] = !f[663] && f[453] && f[303] && f[150]; // c0t290i29
	assign leaf[462] = f[663] && !f[498] && !f[630] && !f[689]; // c0t290i29
	assign leaf[463] = f[663] && !f[498] && !f[630] && f[689]; // c0t290i29
	assign leaf[464] = f[663] && !f[498] && f[630] && !f[604]; // c0t290i29
	assign leaf[465] = f[663] && !f[498] && f[630] && f[604]; // c0t290i29
	assign leaf[466] = f[663] && f[498] && !f[347] && !f[214]; // c0t290i29
	assign leaf[467] = f[663] && f[498] && !f[347] && f[214]; // c0t290i29
	assign leaf[468] = f[663] && f[498] && f[347] && !f[600]; // c0t290i29
	assign leaf[469] = f[663] && f[498] && f[347] && f[600]; // c0t290i29
	assign leaf[470] = !f[444] && !f[213] && !f[240] && !f[326]; // c0t300i30
	assign leaf[471] = !f[444] && !f[213] && !f[240] && f[326]; // c0t300i30
	assign leaf[472] = !f[444] && !f[213] && f[240] && !f[542]; // c0t300i30
	assign leaf[473] = !f[444] && !f[213] && f[240] && f[542]; // c0t300i30
	assign leaf[474] = !f[444] && f[213] && !f[516] && !f[378]; // c0t300i30
	assign leaf[475] = !f[444] && f[213] && !f[516] && f[378]; // c0t300i30
	assign leaf[476] = !f[444] && f[213] && f[516] && !f[658]; // c0t300i30
	assign leaf[477] = !f[444] && f[213] && f[516] && f[658]; // c0t300i30
	assign leaf[478] = f[444] && !f[152] && !f[437] && !f[601]; // c0t300i30
	assign leaf[479] = f[444] && !f[152] && !f[437] && f[601]; // c0t300i30
	assign leaf[480] = f[444] && !f[152] && f[437]; // c0t300i30
	assign leaf[481] = f[444] && f[152] && !f[302] && !f[299]; // c0t300i30
	assign leaf[482] = f[444] && f[152] && !f[302] && f[299]; // c0t300i30
	assign leaf[483] = f[444] && f[152] && f[302]; // c0t300i30
	assign leaf[484] = !f[204] && !f[664] && !f[415] && !f[241]; // c0t310i31
	assign leaf[485] = !f[204] && !f[664] && !f[415] && f[241]; // c0t310i31
	assign leaf[486] = !f[204] && !f[664] && f[415] && !f[436]; // c0t310i31
	assign leaf[487] = !f[204] && !f[664] && f[415] && f[436]; // c0t310i31
	assign leaf[488] = !f[204] && f[664] && !f[269]; // c0t310i31
	assign leaf[489] = !f[204] && f[664] && f[269]; // c0t310i31
	assign leaf[490] = f[204] && !f[398] && !f[399] && !f[272]; // c0t310i31
	assign leaf[491] = f[204] && !f[398] && !f[399] && f[272]; // c0t310i31
	assign leaf[492] = f[204] && !f[398] && f[399] && !f[513]; // c0t310i31
	assign leaf[493] = f[204] && !f[398] && f[399] && f[513]; // c0t310i31
	assign leaf[494] = f[204] && f[398] && !f[470] && !f[629]; // c0t310i31
	assign leaf[495] = f[204] && f[398] && !f[470] && f[629]; // c0t310i31
	assign leaf[496] = f[204] && f[398] && f[470] && !f[378]; // c0t310i31
	assign leaf[497] = f[204] && f[398] && f[470] && f[378]; // c0t310i31
	assign leaf[498] = !f[688] && !f[103] && !f[663] && !f[406]; // c0t320i32
	assign leaf[499] = !f[688] && !f[103] && !f[663] && f[406]; // c0t320i32
	assign leaf[500] = !f[688] && !f[103] && f[663] && !f[659]; // c0t320i32
	assign leaf[501] = !f[688] && !f[103] && f[663] && f[659]; // c0t320i32
	assign leaf[502] = !f[688] && f[103] && !f[517] && !f[301]; // c0t320i32
	assign leaf[503] = !f[688] && f[103] && !f[517] && f[301]; // c0t320i32
	assign leaf[504] = !f[688] && f[103] && f[517] && !f[604]; // c0t320i32
	assign leaf[505] = !f[688] && f[103] && f[517] && f[604]; // c0t320i32
	assign leaf[506] = f[688] && !f[657] && !f[574] && !f[156]; // c0t320i32
	assign leaf[507] = f[688] && !f[657] && !f[574] && f[156]; // c0t320i32
	assign leaf[508] = f[688] && !f[657] && f[574]; // c0t320i32
	assign leaf[509] = f[688] && f[657] && !f[571] && !f[347]; // c0t320i32
	assign leaf[510] = f[688] && f[657] && !f[571] && f[347]; // c0t320i32
	assign leaf[511] = f[688] && f[657] && f[571] && !f[523]; // c0t320i32
	assign leaf[512] = f[688] && f[657] && f[571] && f[523]; // c0t320i32
	assign leaf[513] = !f[571] && !f[436] && !f[360] && !f[512]; // c0t330i33
	assign leaf[514] = !f[571] && !f[436] && !f[360] && f[512]; // c0t330i33
	assign leaf[515] = !f[571] && !f[436] && f[360] && !f[275]; // c0t330i33
	assign leaf[516] = !f[571] && !f[436] && f[360] && f[275]; // c0t330i33
	assign leaf[517] = !f[571] && f[436] && !f[569] && !f[331]; // c0t330i33
	assign leaf[518] = !f[571] && f[436] && !f[569] && f[331]; // c0t330i33
	assign leaf[519] = !f[571] && f[436] && f[569] && !f[461]; // c0t330i33
	assign leaf[520] = !f[571] && f[436] && f[569] && f[461]; // c0t330i33
	assign leaf[521] = f[571] && !f[597] && !f[269] && !f[436]; // c0t330i33
	assign leaf[522] = f[571] && !f[597] && !f[269] && f[436]; // c0t330i33
	assign leaf[523] = f[571] && !f[597] && f[269] && !f[187]; // c0t330i33
	assign leaf[524] = f[571] && !f[597] && f[269] && f[187]; // c0t330i33
	assign leaf[525] = f[571] && f[597] && !f[608] && !f[300]; // c0t330i33
	assign leaf[526] = f[571] && f[597] && !f[608] && f[300]; // c0t330i33
	assign leaf[527] = f[571] && f[597] && f[608] && !f[498]; // c0t330i33
	assign leaf[528] = f[571] && f[597] && f[608] && f[498]; // c0t330i33
	assign leaf[529] = !f[514] && !f[510] && !f[512] && !f[508]; // c0t340i34
	assign leaf[530] = !f[514] && !f[510] && !f[512] && f[508]; // c0t340i34
	assign leaf[531] = !f[514] && !f[510] && f[512] && !f[323]; // c0t340i34
	assign leaf[532] = !f[514] && !f[510] && f[512] && f[323]; // c0t340i34
	assign leaf[533] = !f[514] && f[510] && !f[246] && !f[272]; // c0t340i34
	assign leaf[534] = !f[514] && f[510] && !f[246] && f[272]; // c0t340i34
	assign leaf[535] = !f[514] && f[510] && f[246] && !f[379]; // c0t340i34
	assign leaf[536] = !f[514] && f[510] && f[246] && f[379]; // c0t340i34
	assign leaf[537] = f[514] && !f[656] && !f[359] && !f[520]; // c0t340i34
	assign leaf[538] = f[514] && !f[656] && !f[359] && f[520]; // c0t340i34
	assign leaf[539] = f[514] && !f[656] && f[359] && !f[398]; // c0t340i34
	assign leaf[540] = f[514] && !f[656] && f[359] && f[398]; // c0t340i34
	assign leaf[541] = f[514] && f[656] && !f[521] && !f[153]; // c0t340i34
	assign leaf[542] = f[514] && f[656] && !f[521] && f[153]; // c0t340i34
	assign leaf[543] = f[514] && f[656] && f[521] && !f[483]; // c0t340i34
	assign leaf[544] = f[514] && f[656] && f[521] && f[483]; // c0t340i34
	assign leaf[545] = !f[240] && !f[377] && !f[436] && !f[321]; // c0t350i35
	assign leaf[546] = !f[240] && !f[377] && !f[436] && f[321]; // c0t350i35
	assign leaf[547] = !f[240] && !f[377] && f[436] && !f[270]; // c0t350i35
	assign leaf[548] = !f[240] && !f[377] && f[436] && f[270]; // c0t350i35
	assign leaf[549] = !f[240] && f[377] && !f[461] && !f[218]; // c0t350i35
	assign leaf[550] = !f[240] && f[377] && !f[461] && f[218]; // c0t350i35
	assign leaf[551] = !f[240] && f[377] && f[461] && !f[380]; // c0t350i35
	assign leaf[552] = !f[240] && f[377] && f[461] && f[380]; // c0t350i35
	assign leaf[553] = f[240] && !f[297] && !f[271] && !f[275]; // c0t350i35
	assign leaf[554] = f[240] && !f[297] && !f[271] && f[275]; // c0t350i35
	assign leaf[555] = f[240] && !f[297] && f[271] && !f[321]; // c0t350i35
	assign leaf[556] = f[240] && !f[297] && f[271] && f[321]; // c0t350i35
	assign leaf[557] = f[240] && f[297] && !f[486] && !f[606]; // c0t350i35
	assign leaf[558] = f[240] && f[297] && !f[486] && f[606]; // c0t350i35
	assign leaf[559] = f[240] && f[297] && f[486] && !f[375]; // c0t350i35
	assign leaf[560] = f[240] && f[297] && f[486] && f[375]; // c0t350i35
	assign leaf[561] = !f[711] && !f[609] && !f[177] && !f[415]; // c0t360i36
	assign leaf[562] = !f[711] && !f[609] && !f[177] && f[415]; // c0t360i36
	assign leaf[563] = !f[711] && !f[609] && f[177] && !f[572]; // c0t360i36
	assign leaf[564] = !f[711] && !f[609] && f[177] && f[572]; // c0t360i36
	assign leaf[565] = !f[711] && f[609] && !f[471] && !f[662]; // c0t360i36
	assign leaf[566] = !f[711] && f[609] && !f[471] && f[662]; // c0t360i36
	assign leaf[567] = !f[711] && f[609] && f[471] && !f[346]; // c0t360i36
	assign leaf[568] = !f[711] && f[609] && f[471] && f[346]; // c0t360i36
	assign leaf[569] = f[711] && !f[573]; // c0t360i36
	assign leaf[570] = f[711] && f[573]; // c0t360i36
	assign leaf[571] = !f[213] && !f[408] && !f[377] && !f[461]; // c0t370i37
	assign leaf[572] = !f[213] && !f[408] && !f[377] && f[461]; // c0t370i37
	assign leaf[573] = !f[213] && !f[408] && f[377] && !f[437]; // c0t370i37
	assign leaf[574] = !f[213] && !f[408] && f[377] && f[437]; // c0t370i37
	assign leaf[575] = !f[213] && f[408] && !f[268] && !f[151]; // c0t370i37
	assign leaf[576] = !f[213] && f[408] && !f[268] && f[151]; // c0t370i37
	assign leaf[577] = !f[213] && f[408] && f[268] && !f[490]; // c0t370i37
	assign leaf[578] = !f[213] && f[408] && f[268] && f[490]; // c0t370i37
	assign leaf[579] = f[213] && !f[711] && !f[634] && !f[580]; // c0t370i37
	assign leaf[580] = f[213] && !f[711] && !f[634] && f[580]; // c0t370i37
	assign leaf[581] = f[213] && !f[711] && f[634] && !f[466]; // c0t370i37
	assign leaf[582] = f[213] && !f[711] && f[634] && f[466]; // c0t370i37
	assign leaf[583] = f[213] && f[711] && !f[295]; // c0t370i37
	assign leaf[584] = f[213] && f[711] && f[295]; // c0t370i37
	assign leaf[585] = !f[378] && !f[517] && !f[629] && !f[684]; // c0t380i38
	assign leaf[586] = !f[378] && !f[517] && !f[629] && f[684]; // c0t380i38
	assign leaf[587] = !f[378] && !f[517] && f[629] && !f[323]; // c0t380i38
	assign leaf[588] = !f[378] && !f[517] && f[629] && f[323]; // c0t380i38
	assign leaf[589] = !f[378] && f[517] && !f[427] && !f[377]; // c0t380i38
	assign leaf[590] = !f[378] && f[517] && !f[427] && f[377]; // c0t380i38
	assign leaf[591] = !f[378] && f[517] && f[427] && !f[330]; // c0t380i38
	assign leaf[592] = !f[378] && f[517] && f[427] && f[330]; // c0t380i38
	assign leaf[593] = f[378] && !f[216] && !f[376] && !f[606]; // c0t380i38
	assign leaf[594] = f[378] && !f[216] && !f[376] && f[606]; // c0t380i38
	assign leaf[595] = f[378] && !f[216] && f[376] && !f[406]; // c0t380i38
	assign leaf[596] = f[378] && !f[216] && f[376] && f[406]; // c0t380i38
	assign leaf[597] = f[378] && f[216] && !f[568] && !f[570]; // c0t380i38
	assign leaf[598] = f[378] && f[216] && !f[568] && f[570]; // c0t380i38
	assign leaf[599] = f[378] && f[216] && f[568] && !f[326]; // c0t380i38
	assign leaf[600] = f[378] && f[216] && f[568] && f[326]; // c0t380i38
	assign leaf[601] = !f[240] && !f[326] && !f[436] && !f[128]; // c0t390i39
	assign leaf[602] = !f[240] && !f[326] && !f[436] && f[128]; // c0t390i39
	assign leaf[603] = !f[240] && !f[326] && f[436] && !f[218]; // c0t390i39
	assign leaf[604] = !f[240] && !f[326] && f[436] && f[218]; // c0t390i39
	assign leaf[605] = !f[240] && f[326] && !f[236] && !f[381]; // c0t390i39
	assign leaf[606] = !f[240] && f[326] && !f[236] && f[381]; // c0t390i39
	assign leaf[607] = !f[240] && f[326] && f[236] && !f[397]; // c0t390i39
	assign leaf[608] = !f[240] && f[326] && f[236] && f[397]; // c0t390i39
	assign leaf[609] = f[240] && !f[326] && !f[538] && !f[466]; // c0t390i39
	assign leaf[610] = f[240] && !f[326] && !f[538] && f[466]; // c0t390i39
	assign leaf[611] = f[240] && !f[326] && f[538] && !f[608]; // c0t390i39
	assign leaf[612] = f[240] && !f[326] && f[538] && f[608]; // c0t390i39
	assign leaf[613] = f[240] && f[326] && !f[298] && !f[355]; // c0t390i39
	assign leaf[614] = f[240] && f[326] && !f[298] && f[355]; // c0t390i39
	assign leaf[615] = f[240] && f[326] && f[298] && !f[354]; // c0t390i39
	assign leaf[616] = f[240] && f[326] && f[298] && f[354]; // c0t390i39
	assign leaf[617] = !f[688] && !f[453] && !f[298] && !f[300]; // c0t400i40
	assign leaf[618] = !f[688] && !f[453] && !f[298] && f[300]; // c0t400i40
	assign leaf[619] = !f[688] && !f[453] && f[298] && !f[459]; // c0t400i40
	assign leaf[620] = !f[688] && !f[453] && f[298] && f[459]; // c0t400i40
	assign leaf[621] = !f[688] && f[453] && !f[459] && !f[383]; // c0t400i40
	assign leaf[622] = !f[688] && f[453] && !f[459] && f[383]; // c0t400i40
	assign leaf[623] = !f[688] && f[453] && f[459] && !f[572]; // c0t400i40
	assign leaf[624] = !f[688] && f[453] && f[459] && f[572]; // c0t400i40
	assign leaf[625] = f[688] && !f[657] && !f[549]; // c0t400i40
	assign leaf[626] = f[688] && !f[657] && f[549] && !f[273]; // c0t400i40
	assign leaf[627] = f[688] && !f[657] && f[549] && f[273]; // c0t400i40
	assign leaf[628] = f[688] && f[657] && !f[186] && !f[655]; // c0t400i40
	assign leaf[629] = f[688] && f[657] && !f[186] && f[655]; // c0t400i40
	assign leaf[630] = f[688] && f[657] && f[186] && !f[272]; // c0t400i40
	assign leaf[631] = f[688] && f[657] && f[186] && f[272]; // c0t400i40
	assign leaf[632] = !f[444] && !f[319] && !f[494] && !f[413]; // c0t410i41
	assign leaf[633] = !f[444] && !f[319] && !f[494] && f[413]; // c0t410i41
	assign leaf[634] = !f[444] && !f[319] && f[494] && !f[657]; // c0t410i41
	assign leaf[635] = !f[444] && !f[319] && f[494] && f[657]; // c0t410i41
	assign leaf[636] = !f[444] && f[319] && !f[605] && !f[493]; // c0t410i41
	assign leaf[637] = !f[444] && f[319] && !f[605] && f[493]; // c0t410i41
	assign leaf[638] = !f[444] && f[319] && f[605] && !f[320]; // c0t410i41
	assign leaf[639] = !f[444] && f[319] && f[605] && f[320]; // c0t410i41
	assign leaf[640] = f[444] && !f[152] && !f[289]; // c0t410i41
	assign leaf[641] = f[444] && !f[152] && f[289] && !f[600]; // c0t410i41
	assign leaf[642] = f[444] && !f[152] && f[289] && f[600]; // c0t410i41
	assign leaf[643] = f[444] && f[152] && !f[483]; // c0t410i41
	assign leaf[644] = f[444] && f[152] && f[483] && !f[302]; // c0t410i41
	assign leaf[645] = f[444] && f[152] && f[483] && f[302]; // c0t410i41
	assign leaf[646] = !f[347] && !f[466] && !f[404] && !f[293]; // c0t420i42
	assign leaf[647] = !f[347] && !f[466] && !f[404] && f[293]; // c0t420i42
	assign leaf[648] = !f[347] && !f[466] && f[404] && !f[465]; // c0t420i42
	assign leaf[649] = !f[347] && !f[466] && f[404] && f[465]; // c0t420i42
	assign leaf[650] = !f[347] && f[466] && !f[127] && !f[329]; // c0t420i42
	assign leaf[651] = !f[347] && f[466] && !f[127] && f[329]; // c0t420i42
	assign leaf[652] = !f[347] && f[466] && f[127] && !f[344]; // c0t420i42
	assign leaf[653] = !f[347] && f[466] && f[127] && f[344]; // c0t420i42
	assign leaf[654] = f[347] && !f[493] && !f[348] && !f[551]; // c0t420i42
	assign leaf[655] = f[347] && !f[493] && !f[348] && f[551]; // c0t420i42
	assign leaf[656] = f[347] && !f[493] && f[348] && !f[273]; // c0t420i42
	assign leaf[657] = f[347] && !f[493] && f[348] && f[273]; // c0t420i42
	assign leaf[658] = f[347] && f[493] && !f[577] && !f[523]; // c0t420i42
	assign leaf[659] = f[347] && f[493] && !f[577] && f[523]; // c0t420i42
	assign leaf[660] = f[347] && f[493] && f[577] && !f[491]; // c0t420i42
	assign leaf[661] = f[347] && f[493] && f[577] && f[491]; // c0t420i42
	assign leaf[662] = !f[408] && !f[491] && !f[209] && !f[150]; // c0t430i43
	assign leaf[663] = !f[408] && !f[491] && !f[209] && f[150]; // c0t430i43
	assign leaf[664] = !f[408] && !f[491] && f[209] && !f[488]; // c0t430i43
	assign leaf[665] = !f[408] && !f[491] && f[209] && f[488]; // c0t430i43
	assign leaf[666] = !f[408] && f[491] && !f[210] && !f[576]; // c0t430i43
	assign leaf[667] = !f[408] && f[491] && !f[210] && f[576]; // c0t430i43
	assign leaf[668] = !f[408] && f[491] && f[210] && !f[410]; // c0t430i43
	assign leaf[669] = !f[408] && f[491] && f[210] && f[410]; // c0t430i43
	assign leaf[670] = f[408] && !f[268] && !f[427]; // c0t430i43
	assign leaf[671] = f[408] && !f[268] && f[427] && !f[595]; // c0t430i43
	assign leaf[672] = f[408] && !f[268] && f[427] && f[595]; // c0t430i43
	assign leaf[673] = f[408] && f[268] && !f[514] && !f[271]; // c0t430i43
	assign leaf[674] = f[408] && f[268] && !f[514] && f[271]; // c0t430i43
	assign leaf[675] = f[408] && f[268] && f[514] && !f[656]; // c0t430i43
	assign leaf[676] = f[408] && f[268] && f[514] && f[656]; // c0t430i43
	assign leaf[677] = !f[319] && !f[494] && !f[374] && !f[627]; // c0t440i44
	assign leaf[678] = !f[319] && !f[494] && !f[374] && f[627]; // c0t440i44
	assign leaf[679] = !f[319] && !f[494] && f[374] && !f[376]; // c0t440i44
	assign leaf[680] = !f[319] && !f[494] && f[374] && f[376]; // c0t440i44
	assign leaf[681] = !f[319] && f[494] && !f[237] && !f[176]; // c0t440i44
	assign leaf[682] = !f[319] && f[494] && !f[237] && f[176]; // c0t440i44
	assign leaf[683] = !f[319] && f[494] && f[237] && !f[370]; // c0t440i44
	assign leaf[684] = !f[319] && f[494] && f[237] && f[370]; // c0t440i44
	assign leaf[685] = f[319] && !f[543] && !f[233] && !f[409]; // c0t440i44
	assign leaf[686] = f[319] && !f[543] && !f[233] && f[409]; // c0t440i44
	assign leaf[687] = f[319] && !f[543] && f[233] && !f[297]; // c0t440i44
	assign leaf[688] = f[319] && !f[543] && f[233] && f[297]; // c0t440i44
	assign leaf[689] = f[319] && f[543] && !f[541] && !f[625]; // c0t440i44
	assign leaf[690] = f[319] && f[543] && !f[541] && f[625]; // c0t440i44
	assign leaf[691] = f[319] && f[543] && f[541] && !f[160]; // c0t440i44
	assign leaf[692] = f[319] && f[543] && f[541] && f[160]; // c0t440i44
	assign leaf[693] = !f[444] && !f[375] && !f[520] && !f[293]; // c0t450i45
	assign leaf[694] = !f[444] && !f[375] && !f[520] && f[293]; // c0t450i45
	assign leaf[695] = !f[444] && !f[375] && f[520] && !f[373]; // c0t450i45
	assign leaf[696] = !f[444] && !f[375] && f[520] && f[373]; // c0t450i45
	assign leaf[697] = !f[444] && f[375] && !f[486] && !f[352]; // c0t450i45
	assign leaf[698] = !f[444] && f[375] && !f[486] && f[352]; // c0t450i45
	assign leaf[699] = !f[444] && f[375] && f[486] && !f[99]; // c0t450i45
	assign leaf[700] = !f[444] && f[375] && f[486] && f[99]; // c0t450i45
	assign leaf[701] = f[444] && !f[437] && !f[370]; // c0t450i45
	assign leaf[702] = f[444] && !f[437] && f[370] && !f[379]; // c0t450i45
	assign leaf[703] = f[444] && !f[437] && f[370] && f[379]; // c0t450i45
	assign leaf[704] = f[444] && f[437]; // c0t450i45
	assign leaf[705] = !f[434] && !f[664] && !f[379] && !f[332]; // c0t460i46
	assign leaf[706] = !f[434] && !f[664] && !f[379] && f[332]; // c0t460i46
	assign leaf[707] = !f[434] && !f[664] && f[379] && !f[488]; // c0t460i46
	assign leaf[708] = !f[434] && !f[664] && f[379] && f[488]; // c0t460i46
	assign leaf[709] = !f[434] && f[664] && !f[178]; // c0t460i46
	assign leaf[710] = !f[434] && f[664] && f[178] && !f[498]; // c0t460i46
	assign leaf[711] = !f[434] && f[664] && f[178] && f[498]; // c0t460i46
	assign leaf[712] = f[434] && !f[436] && !f[185]; // c0t460i46
	assign leaf[713] = f[434] && !f[436] && f[185] && !f[457]; // c0t460i46
	assign leaf[714] = f[434] && !f[436] && f[185] && f[457]; // c0t460i46
	assign leaf[715] = f[434] && f[436] && !f[433] && !f[595]; // c0t460i46
	assign leaf[716] = f[434] && f[436] && !f[433] && f[595]; // c0t460i46
	assign leaf[717] = f[434] && f[436] && f[433] && !f[414]; // c0t460i46
	assign leaf[718] = f[434] && f[436] && f[433] && f[414]; // c0t460i46
	assign leaf[719] = !f[714] && !f[710] && !f[427] && !f[431]; // c0t470i47
	assign leaf[720] = !f[714] && !f[710] && !f[427] && f[431]; // c0t470i47
	assign leaf[721] = !f[714] && !f[710] && f[427] && !f[377]; // c0t470i47
	assign leaf[722] = !f[714] && !f[710] && f[427] && f[377]; // c0t470i47
	assign leaf[723] = !f[714] && f[710]; // c0t470i47
	assign leaf[724] = f[714] && !f[576]; // c0t470i47
	assign leaf[725] = f[714] && f[576]; // c0t470i47
	assign leaf[726] = !f[238] && !f[219] && !f[266] && !f[464]; // c0t480i48
	assign leaf[727] = !f[238] && !f[219] && !f[266] && f[464]; // c0t480i48
	assign leaf[728] = !f[238] && !f[219] && f[266] && !f[602]; // c0t480i48
	assign leaf[729] = !f[238] && !f[219] && f[266] && f[602]; // c0t480i48
	assign leaf[730] = !f[238] && f[219] && !f[510] && !f[189]; // c0t480i48
	assign leaf[731] = !f[238] && f[219] && !f[510] && f[189]; // c0t480i48
	assign leaf[732] = !f[238] && f[219] && f[510] && !f[241]; // c0t480i48
	assign leaf[733] = !f[238] && f[219] && f[510] && f[241]; // c0t480i48
	assign leaf[734] = f[238] && !f[269] && !f[625] && !f[386]; // c0t480i48
	assign leaf[735] = f[238] && !f[269] && !f[625] && f[386]; // c0t480i48
	assign leaf[736] = f[238] && !f[269] && f[625] && !f[325]; // c0t480i48
	assign leaf[737] = f[238] && !f[269] && f[625] && f[325]; // c0t480i48
	assign leaf[738] = f[238] && f[269] && !f[244] && !f[515]; // c0t480i48
	assign leaf[739] = f[238] && f[269] && !f[244] && f[515]; // c0t480i48
	assign leaf[740] = f[238] && f[269] && f[244] && !f[295]; // c0t480i48
	assign leaf[741] = f[238] && f[269] && f[244] && f[295]; // c0t480i48
	assign leaf[742] = !f[414] && !f[382] && !f[516] && !f[655]; // c0t490i49
	assign leaf[743] = !f[414] && !f[382] && !f[516] && f[655]; // c0t490i49
	assign leaf[744] = !f[414] && !f[382] && f[516] && !f[151]; // c0t490i49
	assign leaf[745] = !f[414] && !f[382] && f[516] && f[151]; // c0t490i49
	assign leaf[746] = !f[414] && f[382] && !f[403] && !f[373]; // c0t490i49
	assign leaf[747] = !f[414] && f[382] && !f[403] && f[373]; // c0t490i49
	assign leaf[748] = !f[414] && f[382] && f[403] && !f[380]; // c0t490i49
	assign leaf[749] = !f[414] && f[382] && f[403] && f[380]; // c0t490i49
	assign leaf[750] = f[414] && !f[190] && !f[329] && !f[273]; // c0t490i49
	assign leaf[751] = f[414] && !f[190] && !f[329] && f[273]; // c0t490i49
	assign leaf[752] = f[414] && !f[190] && f[329] && !f[513]; // c0t490i49
	assign leaf[753] = f[414] && !f[190] && f[329] && f[513]; // c0t490i49
	assign leaf[754] = f[414] && f[190] && !f[521]; // c0t490i49
	assign leaf[755] = f[414] && f[190] && f[521] && !f[492]; // c0t490i49
	assign leaf[756] = f[414] && f[190] && f[521] && f[492]; // c0t490i49
	assign leaf[757] = !f[572] && !f[460] && !f[404] && !f[537]; // c0t500i50
	assign leaf[758] = !f[572] && !f[460] && !f[404] && f[537]; // c0t500i50
	assign leaf[759] = !f[572] && !f[460] && f[404] && !f[266]; // c0t500i50
	assign leaf[760] = !f[572] && !f[460] && f[404] && f[266]; // c0t500i50
	assign leaf[761] = !f[572] && f[460] && !f[570] && !f[189]; // c0t500i50
	assign leaf[762] = !f[572] && f[460] && !f[570] && f[189]; // c0t500i50
	assign leaf[763] = !f[572] && f[460] && f[570] && !f[628]; // c0t500i50
	assign leaf[764] = !f[572] && f[460] && f[570] && f[628]; // c0t500i50
	assign leaf[765] = f[572] && !f[683] && !f[596] && !f[241]; // c0t500i50
	assign leaf[766] = f[572] && !f[683] && !f[596] && f[241]; // c0t500i50
	assign leaf[767] = f[572] && !f[683] && f[596] && !f[245]; // c0t500i50
	assign leaf[768] = f[572] && !f[683] && f[596] && f[245]; // c0t500i50
	assign leaf[769] = f[572] && f[683] && !f[577]; // c0t500i50
	assign leaf[770] = f[572] && f[683] && f[577]; // c0t500i50
	assign leaf[771] = !f[133] && !f[397] && !f[428] && !f[567]; // c0t510i51
	assign leaf[772] = !f[133] && !f[397] && !f[428] && f[567]; // c0t510i51
	assign leaf[773] = !f[133] && !f[397] && f[428] && !f[458]; // c0t510i51
	assign leaf[774] = !f[133] && !f[397] && f[428] && f[458]; // c0t510i51
	assign leaf[775] = !f[133] && f[397] && !f[626] && !f[498]; // c0t510i51
	assign leaf[776] = !f[133] && f[397] && !f[626] && f[498]; // c0t510i51
	assign leaf[777] = !f[133] && f[397] && f[626] && !f[430]; // c0t510i51
	assign leaf[778] = !f[133] && f[397] && f[626] && f[430]; // c0t510i51
	assign leaf[779] = f[133] && !f[653] && !f[516]; // c0t510i51
	assign leaf[780] = f[133] && !f[653] && f[516]; // c0t510i51
	assign leaf[781] = f[133] && f[653] && !f[512]; // c0t510i51
	assign leaf[782] = f[133] && f[653] && f[512]; // c0t510i51
	assign leaf[783] = !f[378] && !f[352] && !f[453] && !f[518]; // c0t520i52
	assign leaf[784] = !f[378] && !f[352] && !f[453] && f[518]; // c0t520i52
	assign leaf[785] = !f[378] && !f[352] && f[453] && !f[661]; // c0t520i52
	assign leaf[786] = !f[378] && !f[352] && f[453] && f[661]; // c0t520i52
	assign leaf[787] = !f[378] && f[352] && !f[431] && !f[320]; // c0t520i52
	assign leaf[788] = !f[378] && f[352] && !f[431] && f[320]; // c0t520i52
	assign leaf[789] = !f[378] && f[352] && f[431] && !f[294]; // c0t520i52
	assign leaf[790] = !f[378] && f[352] && f[431] && f[294]; // c0t520i52
	assign leaf[791] = f[378] && !f[488] && !f[352] && !f[329]; // c0t520i52
	assign leaf[792] = f[378] && !f[488] && !f[352] && f[329]; // c0t520i52
	assign leaf[793] = f[378] && !f[488] && f[352] && !f[377]; // c0t520i52
	assign leaf[794] = f[378] && !f[488] && f[352] && f[377]; // c0t520i52
	assign leaf[795] = f[378] && f[488] && !f[686] && !f[542]; // c0t520i52
	assign leaf[796] = f[378] && f[488] && !f[686] && f[542]; // c0t520i52
	assign leaf[797] = f[378] && f[488] && f[686]; // c0t520i52
	assign leaf[798] = !f[713] && !f[605] && !f[406] && !f[637]; // c0t530i53
	assign leaf[799] = !f[713] && !f[605] && !f[406] && f[637]; // c0t530i53
	assign leaf[800] = !f[713] && !f[605] && f[406] && !f[216]; // c0t530i53
	assign leaf[801] = !f[713] && !f[605] && f[406] && f[216]; // c0t530i53
	assign leaf[802] = !f[713] && f[605] && !f[207] && !f[683]; // c0t530i53
	assign leaf[803] = !f[713] && f[605] && !f[207] && f[683]; // c0t530i53
	assign leaf[804] = !f[713] && f[605] && f[207] && !f[624]; // c0t530i53
	assign leaf[805] = !f[713] && f[605] && f[207] && f[624]; // c0t530i53
	assign leaf[806] = f[713] && !f[295]; // c0t530i53
	assign leaf[807] = f[713] && f[295]; // c0t530i53
	assign leaf[808] = !f[713] && !f[710] && !f[427] && !f[344]; // c0t540i54
	assign leaf[809] = !f[713] && !f[710] && !f[427] && f[344]; // c0t540i54
	assign leaf[810] = !f[713] && !f[710] && f[427] && !f[345]; // c0t540i54
	assign leaf[811] = !f[713] && !f[710] && f[427] && f[345]; // c0t540i54
	assign leaf[812] = !f[713] && f[710]; // c0t540i54
	assign leaf[813] = f[713] && !f[376]; // c0t540i54
	assign leaf[814] = f[713] && f[376]; // c0t540i54
	assign leaf[815] = !f[444] && !f[609] && !f[402] && !f[494]; // c0t550i55
	assign leaf[816] = !f[444] && !f[609] && !f[402] && f[494]; // c0t550i55
	assign leaf[817] = !f[444] && !f[609] && f[402] && !f[347]; // c0t550i55
	assign leaf[818] = !f[444] && !f[609] && f[402] && f[347]; // c0t550i55
	assign leaf[819] = !f[444] && f[609] && !f[180] && !f[232]; // c0t550i55
	assign leaf[820] = !f[444] && f[609] && !f[180] && f[232]; // c0t550i55
	assign leaf[821] = !f[444] && f[609] && f[180] && !f[347]; // c0t550i55
	assign leaf[822] = !f[444] && f[609] && f[180] && f[347]; // c0t550i55
	assign leaf[823] = f[444] && !f[152] && !f[317]; // c0t550i55
	assign leaf[824] = f[444] && !f[152] && f[317] && !f[359]; // c0t550i55
	assign leaf[825] = f[444] && !f[152] && f[317] && f[359]; // c0t550i55
	assign leaf[826] = f[444] && f[152] && !f[272]; // c0t550i55
	assign leaf[827] = f[444] && f[152] && f[272]; // c0t550i55
	assign leaf[828] = !f[416] && !f[214] && !f[241] && !f[438]; // c0t560i56
	assign leaf[829] = !f[416] && !f[214] && !f[241] && f[438]; // c0t560i56
	assign leaf[830] = !f[416] && !f[214] && f[241] && !f[542]; // c0t560i56
	assign leaf[831] = !f[416] && !f[214] && f[241] && f[542]; // c0t560i56
	assign leaf[832] = !f[416] && f[214] && !f[516] && !f[380]; // c0t560i56
	assign leaf[833] = !f[416] && f[214] && !f[516] && f[380]; // c0t560i56
	assign leaf[834] = !f[416] && f[214] && f[516] && !f[186]; // c0t560i56
	assign leaf[835] = !f[416] && f[214] && f[516] && f[186]; // c0t560i56
	assign leaf[836] = f[416] && !f[398]; // c0t560i56
	assign leaf[837] = f[416] && f[398] && !f[289]; // c0t560i56
	assign leaf[838] = f[416] && f[398] && f[289] && !f[430]; // c0t560i56
	assign leaf[839] = f[416] && f[398] && f[289] && f[430]; // c0t560i56
	assign leaf[840] = !f[434] && !f[664] && !f[433] && !f[547]; // c0t570i57
	assign leaf[841] = !f[434] && !f[664] && !f[433] && f[547]; // c0t570i57
	assign leaf[842] = !f[434] && !f[664] && f[433] && !f[348]; // c0t570i57
	assign leaf[843] = !f[434] && !f[664] && f[433] && f[348]; // c0t570i57
	assign leaf[844] = !f[434] && f[664] && !f[151]; // c0t570i57
	assign leaf[845] = !f[434] && f[664] && f[151]; // c0t570i57
	assign leaf[846] = f[434] && !f[456] && !f[386]; // c0t570i57
	assign leaf[847] = f[434] && !f[456] && f[386]; // c0t570i57
	assign leaf[848] = f[434] && f[456] && !f[461] && !f[267]; // c0t570i57
	assign leaf[849] = f[434] && f[456] && !f[461] && f[267]; // c0t570i57
	assign leaf[850] = f[434] && f[456] && f[461] && !f[357]; // c0t570i57
	assign leaf[851] = f[434] && f[456] && f[461] && f[357]; // c0t570i57
	assign leaf[852] = !f[688] && !f[663] && !f[712] && !f[397]; // c0t580i58
	assign leaf[853] = !f[688] && !f[663] && !f[712] && f[397]; // c0t580i58
	assign leaf[854] = !f[688] && !f[663] && f[712] && !f[573]; // c0t580i58
	assign leaf[855] = !f[688] && !f[663] && f[712] && f[573]; // c0t580i58
	assign leaf[856] = !f[688] && f[663] && !f[659]; // c0t580i58
	assign leaf[857] = !f[688] && f[663] && f[659]; // c0t580i58
	assign leaf[858] = f[688] && !f[548] && !f[287] && !f[356]; // c0t580i58
	assign leaf[859] = f[688] && !f[548] && !f[287] && f[356]; // c0t580i58
	assign leaf[860] = f[688] && !f[548] && f[287]; // c0t580i58
	assign leaf[861] = f[688] && f[548]; // c0t580i58
	assign leaf[862] = !f[380] && !f[512] && !f[271] && !f[403]; // c0t590i59
	assign leaf[863] = !f[380] && !f[512] && !f[271] && f[403]; // c0t590i59
	assign leaf[864] = !f[380] && !f[512] && f[271] && !f[462]; // c0t590i59
	assign leaf[865] = !f[380] && !f[512] && f[271] && f[462]; // c0t590i59
	assign leaf[866] = !f[380] && f[512] && !f[429] && !f[359]; // c0t590i59
	assign leaf[867] = !f[380] && f[512] && !f[429] && f[359]; // c0t590i59
	assign leaf[868] = !f[380] && f[512] && f[429] && !f[353]; // c0t590i59
	assign leaf[869] = !f[380] && f[512] && f[429] && f[353]; // c0t590i59
	assign leaf[870] = f[380] && !f[268] && !f[314] && !f[126]; // c0t590i59
	assign leaf[871] = f[380] && !f[268] && !f[314] && f[126]; // c0t590i59
	assign leaf[872] = f[380] && !f[268] && f[314]; // c0t590i59
	assign leaf[873] = f[380] && f[268] && !f[325] && !f[329]; // c0t590i59
	assign leaf[874] = f[380] && f[268] && !f[325] && f[329]; // c0t590i59
	assign leaf[875] = f[380] && f[268] && f[325] && !f[596]; // c0t590i59
	assign leaf[876] = f[380] && f[268] && f[325] && f[596]; // c0t590i59
	assign leaf[877] = !f[605] && !f[321] && !f[320] && !f[431]; // c0t600i60
	assign leaf[878] = !f[605] && !f[321] && !f[320] && f[431]; // c0t600i60
	assign leaf[879] = !f[605] && !f[321] && f[320] && !f[468]; // c0t600i60
	assign leaf[880] = !f[605] && !f[321] && f[320] && f[468]; // c0t600i60
	assign leaf[881] = !f[605] && f[321] && !f[153] && !f[480]; // c0t600i60
	assign leaf[882] = !f[605] && f[321] && !f[153] && f[480]; // c0t600i60
	assign leaf[883] = !f[605] && f[321] && f[153] && !f[401]; // c0t600i60
	assign leaf[884] = !f[605] && f[321] && f[153] && f[401]; // c0t600i60
	assign leaf[885] = f[605] && !f[207] && !f[492] && !f[273]; // c0t600i60
	assign leaf[886] = f[605] && !f[207] && !f[492] && f[273]; // c0t600i60
	assign leaf[887] = f[605] && !f[207] && f[492] && !f[128]; // c0t600i60
	assign leaf[888] = f[605] && !f[207] && f[492] && f[128]; // c0t600i60
	assign leaf[889] = f[605] && f[207] && !f[185] && !f[354]; // c0t600i60
	assign leaf[890] = f[605] && f[207] && !f[185] && f[354]; // c0t600i60
	assign leaf[891] = f[605] && f[207] && f[185] && !f[316]; // c0t600i60
	assign leaf[892] = f[605] && f[207] && f[185] && f[316]; // c0t600i60
	assign leaf[893] = !f[572] && !f[547] && !f[376] && !f[460]; // c0t610i61
	assign leaf[894] = !f[572] && !f[547] && !f[376] && f[460]; // c0t610i61
	assign leaf[895] = !f[572] && !f[547] && f[376] && !f[189]; // c0t610i61
	assign leaf[896] = !f[572] && !f[547] && f[376] && f[189]; // c0t610i61
	assign leaf[897] = !f[572] && f[547] && !f[294] && !f[268]; // c0t610i61
	assign leaf[898] = !f[572] && f[547] && !f[294] && f[268]; // c0t610i61
	assign leaf[899] = !f[572] && f[547] && f[294] && !f[576]; // c0t610i61
	assign leaf[900] = !f[572] && f[547] && f[294] && f[576]; // c0t610i61
	assign leaf[901] = f[572] && !f[683] && !f[319] && !f[354]; // c0t610i61
	assign leaf[902] = f[572] && !f[683] && !f[319] && f[354]; // c0t610i61
	assign leaf[903] = f[572] && !f[683] && f[319] && !f[598]; // c0t610i61
	assign leaf[904] = f[572] && !f[683] && f[319] && f[598]; // c0t610i61
	assign leaf[905] = f[572] && f[683]; // c0t610i61
	assign leaf[906] = !f[572] && !f[541] && !f[494] && !f[595]; // c0t620i62
	assign leaf[907] = !f[572] && !f[541] && !f[494] && f[595]; // c0t620i62
	assign leaf[908] = !f[572] && !f[541] && f[494] && !f[316]; // c0t620i62
	assign leaf[909] = !f[572] && !f[541] && f[494] && f[316]; // c0t620i62
	assign leaf[910] = !f[572] && f[541] && !f[353] && !f[485]; // c0t620i62
	assign leaf[911] = !f[572] && f[541] && !f[353] && f[485]; // c0t620i62
	assign leaf[912] = !f[572] && f[541] && f[353] && !f[607]; // c0t620i62
	assign leaf[913] = !f[572] && f[541] && f[353] && f[607]; // c0t620i62
	assign leaf[914] = f[572] && !f[683] && !f[459] && !f[455]; // c0t620i62
	assign leaf[915] = f[572] && !f[683] && !f[459] && f[455]; // c0t620i62
	assign leaf[916] = f[572] && !f[683] && f[459] && !f[686]; // c0t620i62
	assign leaf[917] = f[572] && !f[683] && f[459] && f[686]; // c0t620i62
	assign leaf[918] = f[572] && f[683] && !f[549]; // c0t620i62
	assign leaf[919] = f[572] && f[683] && f[549]; // c0t620i62
	assign leaf[920] = !f[380] && !f[382] && !f[303] && !f[517]; // c0t630i63
	assign leaf[921] = !f[380] && !f[382] && !f[303] && f[517]; // c0t630i63
	assign leaf[922] = !f[380] && !f[382] && f[303] && !f[385]; // c0t630i63
	assign leaf[923] = !f[380] && !f[382] && f[303] && f[385]; // c0t630i63
	assign leaf[924] = !f[380] && f[382] && !f[403] && !f[385]; // c0t630i63
	assign leaf[925] = !f[380] && f[382] && !f[403] && f[385]; // c0t630i63
	assign leaf[926] = !f[380] && f[382] && f[403] && !f[408]; // c0t630i63
	assign leaf[927] = !f[380] && f[382] && f[403] && f[408]; // c0t630i63
	assign leaf[928] = f[380] && !f[406] && !f[656] && !f[155]; // c0t630i63
	assign leaf[929] = f[380] && !f[406] && !f[656] && f[155]; // c0t630i63
	assign leaf[930] = f[380] && !f[406] && f[656] && !f[492]; // c0t630i63
	assign leaf[931] = f[380] && !f[406] && f[656] && f[492]; // c0t630i63
	assign leaf[932] = f[380] && f[406] && !f[244]; // c0t630i63
	assign leaf[933] = f[380] && f[406] && f[244] && !f[129]; // c0t630i63
	assign leaf[934] = f[380] && f[406] && f[244] && f[129]; // c0t630i63
	assign leaf[935] = !f[412] && !f[238] && !f[269] && !f[437]; // c0t640i64
	assign leaf[936] = !f[412] && !f[238] && !f[269] && f[437]; // c0t640i64
	assign leaf[937] = !f[412] && !f[238] && f[269] && !f[354]; // c0t640i64
	assign leaf[938] = !f[412] && !f[238] && f[269] && f[354]; // c0t640i64
	assign leaf[939] = !f[412] && f[238] && !f[331] && !f[216]; // c0t640i64
	assign leaf[940] = !f[412] && f[238] && !f[331] && f[216]; // c0t640i64
	assign leaf[941] = !f[412] && f[238] && f[331] && !f[329]; // c0t640i64
	assign leaf[942] = !f[412] && f[238] && f[331] && f[329]; // c0t640i64
	assign leaf[943] = f[412] && !f[572] && !f[682] && !f[210]; // c0t640i64
	assign leaf[944] = f[412] && !f[572] && !f[682] && f[210]; // c0t640i64
	assign leaf[945] = f[412] && !f[572] && f[682] && !f[652]; // c0t640i64
	assign leaf[946] = f[412] && !f[572] && f[682] && f[652]; // c0t640i64
	assign leaf[947] = f[412] && f[572] && !f[321] && !f[387]; // c0t640i64
	assign leaf[948] = f[412] && f[572] && !f[321] && f[387]; // c0t640i64
	assign leaf[949] = f[412] && f[572] && f[321] && !f[403]; // c0t640i64
	assign leaf[950] = f[412] && f[572] && f[321] && f[403]; // c0t640i64
	assign leaf[951] = !f[602] && !f[456] && !f[461] && !f[427]; // c0t650i65
	assign leaf[952] = !f[602] && !f[456] && !f[461] && f[427]; // c0t650i65
	assign leaf[953] = !f[602] && !f[456] && f[461]; // c0t650i65
	assign leaf[954] = !f[602] && f[456] && !f[462] && !f[409]; // c0t650i65
	assign leaf[955] = !f[602] && f[456] && !f[462] && f[409]; // c0t650i65
	assign leaf[956] = !f[602] && f[456] && f[462] && !f[460]; // c0t650i65
	assign leaf[957] = !f[602] && f[456] && f[462] && f[460]; // c0t650i65
	assign leaf[958] = f[602] && !f[236] && !f[350] && !f[549]; // c0t650i65
	assign leaf[959] = f[602] && !f[236] && !f[350] && f[549]; // c0t650i65
	assign leaf[960] = f[602] && !f[236] && f[350] && !f[189]; // c0t650i65
	assign leaf[961] = f[602] && !f[236] && f[350] && f[189]; // c0t650i65
	assign leaf[962] = f[602] && f[236] && !f[463] && !f[483]; // c0t650i65
	assign leaf[963] = f[602] && f[236] && !f[463] && f[483]; // c0t650i65
	assign leaf[964] = f[602] && f[236] && f[463] && !f[321]; // c0t650i65
	assign leaf[965] = f[602] && f[236] && f[463] && f[321]; // c0t650i65
	assign leaf[966] = !f[572] && !f[684] && !f[541] && !f[629]; // c0t660i66
	assign leaf[967] = !f[572] && !f[684] && !f[541] && f[629]; // c0t660i66
	assign leaf[968] = !f[572] && !f[684] && f[541] && !f[212]; // c0t660i66
	assign leaf[969] = !f[572] && !f[684] && f[541] && f[212]; // c0t660i66
	assign leaf[970] = !f[572] && f[684] && !f[574] && !f[353]; // c0t660i66
	assign leaf[971] = !f[572] && f[684] && !f[574] && f[353]; // c0t660i66
	assign leaf[972] = !f[572] && f[684] && f[574] && !f[596]; // c0t660i66
	assign leaf[973] = !f[572] && f[684] && f[574] && f[596]; // c0t660i66
	assign leaf[974] = f[572] && !f[683] && !f[598] && !f[319]; // c0t660i66
	assign leaf[975] = f[572] && !f[683] && !f[598] && f[319]; // c0t660i66
	assign leaf[976] = f[572] && !f[683] && f[598] && !f[608]; // c0t660i66
	assign leaf[977] = f[572] && !f[683] && f[598] && f[608]; // c0t660i66
	assign leaf[978] = f[572] && f[683] && !f[548]; // c0t660i66
	assign leaf[979] = f[572] && f[683] && f[548]; // c0t660i66
	assign leaf[980] = !f[444] && !f[633] && !f[580] && !f[713]; // c0t670i67
	assign leaf[981] = !f[444] && !f[633] && !f[580] && f[713]; // c0t670i67
	assign leaf[982] = !f[444] && !f[633] && f[580] && !f[354]; // c0t670i67
	assign leaf[983] = !f[444] && !f[633] && f[580] && f[354]; // c0t670i67
	assign leaf[984] = !f[444] && f[633] && !f[552] && !f[658]; // c0t670i67
	assign leaf[985] = !f[444] && f[633] && !f[552] && f[658]; // c0t670i67
	assign leaf[986] = !f[444] && f[633] && f[552] && !f[544]; // c0t670i67
	assign leaf[987] = !f[444] && f[633] && f[552] && f[544]; // c0t670i67
	assign leaf[988] = f[444] && !f[152] && !f[317]; // c0t670i67
	assign leaf[989] = f[444] && !f[152] && f[317]; // c0t670i67
	assign leaf[990] = f[444] && f[152]; // c0t670i67
	assign leaf[991] = !f[444] && !f[516] && !f[379] && !f[486]; // c0t680i68
	assign leaf[992] = !f[444] && !f[516] && !f[379] && f[486]; // c0t680i68
	assign leaf[993] = !f[444] && !f[516] && f[379] && !f[268]; // c0t680i68
	assign leaf[994] = !f[444] && !f[516] && f[379] && f[268]; // c0t680i68
	assign leaf[995] = !f[444] && f[516] && !f[437] && !f[206]; // c0t680i68
	assign leaf[996] = !f[444] && f[516] && !f[437] && f[206]; // c0t680i68
	assign leaf[997] = !f[444] && f[516] && f[437] && !f[596]; // c0t680i68
	assign leaf[998] = !f[444] && f[516] && f[437] && f[596]; // c0t680i68
	assign leaf[999] = f[444] && !f[514] && !f[357]; // c0t680i68
	assign leaf[1000] = f[444] && !f[514] && f[357]; // c0t680i68
	assign leaf[1001] = f[444] && f[514] && !f[602]; // c0t680i68
	assign leaf[1002] = f[444] && f[514] && f[602]; // c0t680i68
	assign leaf[1003] = !f[633] && !f[580] && !f[378] && !f[599]; // c0t690i69
	assign leaf[1004] = !f[633] && !f[580] && !f[378] && f[599]; // c0t690i69
	assign leaf[1005] = !f[633] && !f[580] && f[378] && !f[435]; // c0t690i69
	assign leaf[1006] = !f[633] && !f[580] && f[378] && f[435]; // c0t690i69
	assign leaf[1007] = !f[633] && f[580] && !f[568] && !f[471]; // c0t690i69
	assign leaf[1008] = !f[633] && f[580] && !f[568] && f[471]; // c0t690i69
	assign leaf[1009] = !f[633] && f[580] && f[568] && !f[182]; // c0t690i69
	assign leaf[1010] = !f[633] && f[580] && f[568] && f[182]; // c0t690i69
	assign leaf[1011] = f[633] && !f[234] && !f[205] && !f[686]; // c0t690i69
	assign leaf[1012] = f[633] && !f[234] && !f[205] && f[686]; // c0t690i69
	assign leaf[1013] = f[633] && !f[234] && f[205]; // c0t690i69
	assign leaf[1014] = f[633] && f[234] && !f[629] && !f[179]; // c0t690i69
	assign leaf[1015] = f[633] && f[234] && !f[629] && f[179]; // c0t690i69
	assign leaf[1016] = f[633] && f[234] && f[629] && !f[655]; // c0t690i69
	assign leaf[1017] = f[633] && f[234] && f[629] && f[655]; // c0t690i69
	assign leaf[1018] = !f[380] && !f[456] && !f[424] && !f[267]; // c0t700i70
	assign leaf[1019] = !f[380] && !f[456] && !f[424] && f[267]; // c0t700i70
	assign leaf[1020] = !f[380] && !f[456] && f[424] && !f[439]; // c0t700i70
	assign leaf[1021] = !f[380] && !f[456] && f[424] && f[439]; // c0t700i70
	assign leaf[1022] = !f[380] && f[456] && !f[654] && !f[575]; // c0t700i70
	assign leaf[1023] = !f[380] && f[456] && !f[654] && f[575]; // c0t700i70
	assign leaf[1024] = !f[380] && f[456] && f[654] && !f[512]; // c0t700i70
	assign leaf[1025] = !f[380] && f[456] && f[654] && f[512]; // c0t700i70
	assign leaf[1026] = f[380] && !f[350] && !f[324] && !f[407]; // c0t700i70
	assign leaf[1027] = f[380] && !f[350] && !f[324] && f[407]; // c0t700i70
	assign leaf[1028] = f[380] && !f[350] && f[324] && !f[262]; // c0t700i70
	assign leaf[1029] = f[380] && !f[350] && f[324] && f[262]; // c0t700i70
	assign leaf[1030] = f[380] && f[350] && !f[154] && !f[512]; // c0t700i70
	assign leaf[1031] = f[380] && f[350] && !f[154] && f[512]; // c0t700i70
	assign leaf[1032] = f[380] && f[350] && f[154] && !f[382]; // c0t700i70
	assign leaf[1033] = f[380] && f[350] && f[154] && f[382]; // c0t700i70
	assign leaf[1034] = !f[688] && !f[152] && !f[654] && !f[275]; // c0t710i71
	assign leaf[1035] = !f[688] && !f[152] && !f[654] && f[275]; // c0t710i71
	assign leaf[1036] = !f[688] && !f[152] && f[654] && !f[157]; // c0t710i71
	assign leaf[1037] = !f[688] && !f[152] && f[654] && f[157]; // c0t710i71
	assign leaf[1038] = !f[688] && f[152] && !f[349] && !f[293]; // c0t710i71
	assign leaf[1039] = !f[688] && f[152] && !f[349] && f[293]; // c0t710i71
	assign leaf[1040] = !f[688] && f[152] && f[349] && !f[238]; // c0t710i71
	assign leaf[1041] = !f[688] && f[152] && f[349] && f[238]; // c0t710i71
	assign leaf[1042] = f[688] && !f[657]; // c0t710i71
	assign leaf[1043] = f[688] && f[657] && !f[231]; // c0t710i71
	assign leaf[1044] = f[688] && f[657] && f[231]; // c0t710i71
	assign leaf[1045] = !f[466] && !f[213] && !f[293] && !f[517]; // c0t720i72
	assign leaf[1046] = !f[466] && !f[213] && !f[293] && f[517]; // c0t720i72
	assign leaf[1047] = !f[466] && !f[213] && f[293] && !f[521]; // c0t720i72
	assign leaf[1048] = !f[466] && !f[213] && f[293] && f[521]; // c0t720i72
	assign leaf[1049] = !f[466] && f[213] && !f[513] && !f[410]; // c0t720i72
	assign leaf[1050] = !f[466] && f[213] && !f[513] && f[410]; // c0t720i72
	assign leaf[1051] = !f[466] && f[213] && f[513] && !f[524]; // c0t720i72
	assign leaf[1052] = !f[466] && f[213] && f[513] && f[524]; // c0t720i72
	assign leaf[1053] = f[466] && !f[688] && !f[379] && !f[551]; // c0t720i72
	assign leaf[1054] = f[466] && !f[688] && !f[379] && f[551]; // c0t720i72
	assign leaf[1055] = f[466] && !f[688] && f[379] && !f[659]; // c0t720i72
	assign leaf[1056] = f[466] && !f[688] && f[379] && f[659]; // c0t720i72
	assign leaf[1057] = f[466] && f[688]; // c0t720i72
	assign leaf[1058] = !f[683] && !f[714] && !f[183] && !f[609]; // c0t730i73
	assign leaf[1059] = !f[683] && !f[714] && !f[183] && f[609]; // c0t730i73
	assign leaf[1060] = !f[683] && !f[714] && f[183] && !f[630]; // c0t730i73
	assign leaf[1061] = !f[683] && !f[714] && f[183] && f[630]; // c0t730i73
	assign leaf[1062] = !f[683] && f[714]; // c0t730i73
	assign leaf[1063] = f[683] && !f[185]; // c0t730i73
	assign leaf[1064] = f[683] && f[185] && !f[490] && !f[272]; // c0t730i73
	assign leaf[1065] = f[683] && f[185] && !f[490] && f[272]; // c0t730i73
	assign leaf[1066] = f[683] && f[185] && f[490]; // c0t730i73
	assign leaf[1067] = !f[427] && !f[597] && !f[571] && !f[317]; // c0t740i74
	assign leaf[1068] = !f[427] && !f[597] && !f[571] && f[317]; // c0t740i74
	assign leaf[1069] = !f[427] && !f[597] && f[571] && !f[263]; // c0t740i74
	assign leaf[1070] = !f[427] && !f[597] && f[571] && f[263]; // c0t740i74
	assign leaf[1071] = !f[427] && f[597] && !f[516] && !f[324]; // c0t740i74
	assign leaf[1072] = !f[427] && f[597] && !f[516] && f[324]; // c0t740i74
	assign leaf[1073] = !f[427] && f[597] && f[516] && !f[406]; // c0t740i74
	assign leaf[1074] = !f[427] && f[597] && f[516] && f[406]; // c0t740i74
	assign leaf[1075] = f[427] && !f[569] && !f[431] && !f[324]; // c0t740i74
	assign leaf[1076] = f[427] && !f[569] && !f[431] && f[324]; // c0t740i74
	assign leaf[1077] = f[427] && !f[569] && f[431]; // c0t740i74
	assign leaf[1078] = f[427] && f[569] && !f[458] && !f[548]; // c0t740i74
	assign leaf[1079] = f[427] && f[569] && !f[458] && f[548]; // c0t740i74
	assign leaf[1080] = f[427] && f[569] && f[458] && !f[440]; // c0t740i74
	assign leaf[1081] = f[427] && f[569] && f[458] && f[440]; // c0t740i74
	assign leaf[1082] = !f[602] && !f[576] && !f[460] && !f[205]; // c0t750i75
	assign leaf[1083] = !f[602] && !f[576] && !f[460] && f[205]; // c0t750i75
	assign leaf[1084] = !f[602] && !f[576] && f[460] && !f[351]; // c0t750i75
	assign leaf[1085] = !f[602] && !f[576] && f[460] && f[351]; // c0t750i75
	assign leaf[1086] = !f[602] && f[576] && !f[442] && !f[656]; // c0t750i75
	assign leaf[1087] = !f[602] && f[576] && !f[442] && f[656]; // c0t750i75
	assign leaf[1088] = !f[602] && f[576] && f[442]; // c0t750i75
	assign leaf[1089] = f[602] && !f[323] && !f[600] && !f[626]; // c0t750i75
	assign leaf[1090] = f[602] && !f[323] && !f[600] && f[626]; // c0t750i75
	assign leaf[1091] = f[602] && !f[323] && f[600] && !f[630]; // c0t750i75
	assign leaf[1092] = f[602] && !f[323] && f[600] && f[630]; // c0t750i75
	assign leaf[1093] = f[602] && f[323] && !f[264] && !f[433]; // c0t750i75
	assign leaf[1094] = f[602] && f[323] && !f[264] && f[433]; // c0t750i75
	assign leaf[1095] = f[602] && f[323] && f[264] && !f[626]; // c0t750i75
	assign leaf[1096] = f[602] && f[323] && f[264] && f[626]; // c0t750i75
	assign leaf[1097] = !f[213] && !f[544] && !f[384] && !f[408]; // c0t760i76
	assign leaf[1098] = !f[213] && !f[544] && !f[384] && f[408]; // c0t760i76
	assign leaf[1099] = !f[213] && !f[544] && f[384] && !f[215]; // c0t760i76
	assign leaf[1100] = !f[213] && !f[544] && f[384] && f[215]; // c0t760i76
	assign leaf[1101] = !f[213] && f[544] && !f[296] && !f[481]; // c0t760i76
	assign leaf[1102] = !f[213] && f[544] && !f[296] && f[481]; // c0t760i76
	assign leaf[1103] = !f[213] && f[544] && f[296] && !f[494]; // c0t760i76
	assign leaf[1104] = !f[213] && f[544] && f[296] && f[494]; // c0t760i76
	assign leaf[1105] = f[213] && !f[323] && !f[347] && !f[519]; // c0t760i76
	assign leaf[1106] = f[213] && !f[323] && !f[347] && f[519]; // c0t760i76
	assign leaf[1107] = f[213] && !f[323] && f[347] && !f[316]; // c0t760i76
	assign leaf[1108] = f[213] && !f[323] && f[347] && f[316]; // c0t760i76
	assign leaf[1109] = f[213] && f[323] && !f[153] && !f[428]; // c0t760i76
	assign leaf[1110] = f[213] && f[323] && !f[153] && f[428]; // c0t760i76
	assign leaf[1111] = f[213] && f[323] && f[153] && !f[490]; // c0t760i76
	assign leaf[1112] = f[213] && f[323] && f[153] && f[490]; // c0t760i76
	assign leaf[1113] = !f[434] && !f[486] && !f[489] && !f[276]; // c0t770i77
	assign leaf[1114] = !f[434] && !f[486] && !f[489] && f[276]; // c0t770i77
	assign leaf[1115] = !f[434] && !f[486] && f[489] && !f[354]; // c0t770i77
	assign leaf[1116] = !f[434] && !f[486] && f[489] && f[354]; // c0t770i77
	assign leaf[1117] = !f[434] && f[486] && !f[287] && !f[489]; // c0t770i77
	assign leaf[1118] = !f[434] && f[486] && !f[287] && f[489]; // c0t770i77
	assign leaf[1119] = !f[434] && f[486] && f[287] && !f[291]; // c0t770i77
	assign leaf[1120] = !f[434] && f[486] && f[287] && f[291]; // c0t770i77
	assign leaf[1121] = f[434] && !f[357] && !f[461]; // c0t770i77
	assign leaf[1122] = f[434] && !f[357] && f[461]; // c0t770i77
	assign leaf[1123] = f[434] && f[357] && !f[158] && !f[546]; // c0t770i77
	assign leaf[1124] = f[434] && f[357] && !f[158] && f[546]; // c0t770i77
	assign leaf[1125] = f[434] && f[357] && f[158] && !f[409]; // c0t770i77
	assign leaf[1126] = f[434] && f[357] && f[158] && f[409]; // c0t770i77
	assign leaf[1127] = !f[512] && !f[462] && !f[597] && !f[155]; // c0t780i78
	assign leaf[1128] = !f[512] && !f[462] && !f[597] && f[155]; // c0t780i78
	assign leaf[1129] = !f[512] && !f[462] && f[597] && !f[606]; // c0t780i78
	assign leaf[1130] = !f[512] && !f[462] && f[597] && f[606]; // c0t780i78
	assign leaf[1131] = !f[512] && f[462] && !f[481]; // c0t780i78
	assign leaf[1132] = !f[512] && f[462] && f[481]; // c0t780i78
	assign leaf[1133] = f[512] && !f[654] && !f[575] && !f[484]; // c0t780i78
	assign leaf[1134] = f[512] && !f[654] && !f[575] && f[484]; // c0t780i78
	assign leaf[1135] = f[512] && !f[654] && f[575] && !f[437]; // c0t780i78
	assign leaf[1136] = f[512] && !f[654] && f[575] && f[437]; // c0t780i78
	assign leaf[1137] = f[512] && f[654] && !f[247] && !f[400]; // c0t780i78
	assign leaf[1138] = f[512] && f[654] && !f[247] && f[400]; // c0t780i78
	assign leaf[1139] = f[512] && f[654] && f[247]; // c0t780i78
	assign leaf[1140] = !f[607] && !f[688] && !f[192] && !f[258]; // c0t790i79
	assign leaf[1141] = !f[607] && !f[688] && !f[192] && f[258]; // c0t790i79
	assign leaf[1142] = !f[607] && !f[688] && f[192]; // c0t790i79
	assign leaf[1143] = !f[607] && f[688]; // c0t790i79
	assign leaf[1144] = f[607] && !f[633] && !f[439]; // c0t790i79
	assign leaf[1145] = f[607] && !f[633] && f[439]; // c0t790i79
	assign leaf[1146] = f[607] && f[633] && !f[208] && !f[371]; // c0t790i79
	assign leaf[1147] = f[607] && f[633] && !f[208] && f[371]; // c0t790i79
	assign leaf[1148] = f[607] && f[633] && f[208] && !f[157]; // c0t790i79
	assign leaf[1149] = f[607] && f[633] && f[208] && f[157]; // c0t790i79
	assign leaf[1150] = !f[526] && !f[635] && !f[688] && !f[378]; // c0t800i80
	assign leaf[1151] = !f[526] && !f[635] && !f[688] && f[378]; // c0t800i80
	assign leaf[1152] = !f[526] && !f[635] && f[688]; // c0t800i80
	assign leaf[1153] = !f[526] && f[635] && !f[578]; // c0t800i80
	assign leaf[1154] = !f[526] && f[635] && f[578] && !f[429]; // c0t800i80
	assign leaf[1155] = !f[526] && f[635] && f[578] && f[429]; // c0t800i80
	assign leaf[1156] = f[526] && !f[374] && !f[236] && !f[634]; // c0t800i80
	assign leaf[1157] = f[526] && !f[374] && !f[236] && f[634]; // c0t800i80
	assign leaf[1158] = f[526] && !f[374] && f[236] && !f[179]; // c0t800i80
	assign leaf[1159] = f[526] && !f[374] && f[236] && f[179]; // c0t800i80
	assign leaf[1160] = f[526] && f[374] && !f[544] && !f[233]; // c0t800i80
	assign leaf[1161] = f[526] && f[374] && !f[544] && f[233]; // c0t800i80
	assign leaf[1162] = f[526] && f[374] && f[544]; // c0t800i80
	assign leaf[1163] = !f[386] && !f[497] && !f[354] && !f[511]; // c0t810i81
	assign leaf[1164] = !f[386] && !f[497] && !f[354] && f[511]; // c0t810i81
	assign leaf[1165] = !f[386] && !f[497] && f[354] && !f[509]; // c0t810i81
	assign leaf[1166] = !f[386] && !f[497] && f[354] && f[509]; // c0t810i81
	assign leaf[1167] = !f[386] && f[497] && !f[331] && !f[123]; // c0t810i81
	assign leaf[1168] = !f[386] && f[497] && !f[331] && f[123]; // c0t810i81
	assign leaf[1169] = !f[386] && f[497] && f[331]; // c0t810i81
	assign leaf[1170] = f[386] && !f[410] && !f[387] && !f[466]; // c0t810i81
	assign leaf[1171] = f[386] && !f[410] && !f[387] && f[466]; // c0t810i81
	assign leaf[1172] = f[386] && !f[410] && f[387] && !f[302]; // c0t810i81
	assign leaf[1173] = f[386] && !f[410] && f[387] && f[302]; // c0t810i81
	assign leaf[1174] = f[386] && f[410] && !f[513]; // c0t810i81
	assign leaf[1175] = f[386] && f[410] && f[513] && !f[297]; // c0t810i81
	assign leaf[1176] = f[386] && f[410] && f[513] && f[297]; // c0t810i81
	assign leaf[1177] = !f[434] && !f[459] && !f[349] && !f[547]; // c0t820i82
	assign leaf[1178] = !f[434] && !f[459] && !f[349] && f[547]; // c0t820i82
	assign leaf[1179] = !f[434] && !f[459] && f[349] && !f[426]; // c0t820i82
	assign leaf[1180] = !f[434] && !f[459] && f[349] && f[426]; // c0t820i82
	assign leaf[1181] = !f[434] && f[459] && !f[601] && !f[484]; // c0t820i82
	assign leaf[1182] = !f[434] && f[459] && !f[601] && f[484]; // c0t820i82
	assign leaf[1183] = !f[434] && f[459] && f[601] && !f[656]; // c0t820i82
	assign leaf[1184] = !f[434] && f[459] && f[601] && f[656]; // c0t820i82
	assign leaf[1185] = f[434] && !f[433]; // c0t820i82
	assign leaf[1186] = f[434] && f[433] && !f[431]; // c0t820i82
	assign leaf[1187] = f[434] && f[433] && f[431] && !f[521]; // c0t820i82
	assign leaf[1188] = f[434] && f[433] && f[431] && f[521]; // c0t820i82
	assign leaf[1189] = !f[380] && !f[512] && !f[629] && !f[290]; // c0t830i83
	assign leaf[1190] = !f[380] && !f[512] && !f[629] && f[290]; // c0t830i83
	assign leaf[1191] = !f[380] && !f[512] && f[629] && !f[209]; // c0t830i83
	assign leaf[1192] = !f[380] && !f[512] && f[629] && f[209]; // c0t830i83
	assign leaf[1193] = !f[380] && f[512] && !f[302] && !f[517]; // c0t830i83
	assign leaf[1194] = !f[380] && f[512] && !f[302] && f[517]; // c0t830i83
	assign leaf[1195] = !f[380] && f[512] && f[302] && !f[271]; // c0t830i83
	assign leaf[1196] = !f[380] && f[512] && f[302] && f[271]; // c0t830i83
	assign leaf[1197] = f[380] && !f[297] && !f[184]; // c0t830i83
	assign leaf[1198] = f[380] && !f[297] && f[184]; // c0t830i83
	assign leaf[1199] = f[380] && f[297] && !f[435] && !f[262]; // c0t830i83
	assign leaf[1200] = f[380] && f[297] && !f[435] && f[262]; // c0t830i83
	assign leaf[1201] = f[380] && f[297] && f[435] && !f[406]; // c0t830i83
	assign leaf[1202] = f[380] && f[297] && f[435] && f[406]; // c0t830i83
	assign leaf[1203] = !f[152] && !f[294] && !f[155] && !f[488]; // c0t840i84
	assign leaf[1204] = !f[152] && !f[294] && !f[155] && f[488]; // c0t840i84
	assign leaf[1205] = !f[152] && !f[294] && f[155] && !f[463]; // c0t840i84
	assign leaf[1206] = !f[152] && !f[294] && f[155] && f[463]; // c0t840i84
	assign leaf[1207] = !f[152] && f[294] && !f[100] && !f[351]; // c0t840i84
	assign leaf[1208] = !f[152] && f[294] && !f[100] && f[351]; // c0t840i84
	assign leaf[1209] = !f[152] && f[294] && f[100]; // c0t840i84
	assign leaf[1210] = f[152] && !f[371] && !f[539] && !f[156]; // c0t840i84
	assign leaf[1211] = f[152] && !f[371] && !f[539] && f[156]; // c0t840i84
	assign leaf[1212] = f[152] && !f[371] && f[539] && !f[465]; // c0t840i84
	assign leaf[1213] = f[152] && !f[371] && f[539] && f[465]; // c0t840i84
	assign leaf[1214] = f[152] && f[371] && !f[455]; // c0t840i84
	assign leaf[1215] = f[152] && f[371] && f[455] && !f[214]; // c0t840i84
	assign leaf[1216] = f[152] && f[371] && f[455] && f[214]; // c0t840i84
	assign leaf[1217] = !f[681] && !f[345] && !f[375] && !f[498]; // c0t850i85
	assign leaf[1218] = !f[681] && !f[345] && !f[375] && f[498]; // c0t850i85
	assign leaf[1219] = !f[681] && !f[345] && f[375] && !f[429]; // c0t850i85
	assign leaf[1220] = !f[681] && !f[345] && f[375] && f[429]; // c0t850i85
	assign leaf[1221] = !f[681] && f[345] && !f[376] && !f[570]; // c0t850i85
	assign leaf[1222] = !f[681] && f[345] && !f[376] && f[570]; // c0t850i85
	assign leaf[1223] = !f[681] && f[345] && f[376] && !f[264]; // c0t850i85
	assign leaf[1224] = !f[681] && f[345] && f[376] && f[264]; // c0t850i85
	assign leaf[1225] = f[681] && !f[599] && !f[354] && !f[523]; // c0t850i85
	assign leaf[1226] = f[681] && !f[599] && !f[354] && f[523]; // c0t850i85
	assign leaf[1227] = f[681] && !f[599] && f[354]; // c0t850i85
	assign leaf[1228] = f[681] && f[599] && !f[575]; // c0t850i85
	assign leaf[1229] = f[681] && f[599] && f[575]; // c0t850i85
	assign leaf[1230] = !f[633] && !f[683] && !f[608] && !f[378]; // c0t860i86
	assign leaf[1231] = !f[633] && !f[683] && !f[608] && f[378]; // c0t860i86
	assign leaf[1232] = !f[633] && !f[683] && f[608]; // c0t860i86
	assign leaf[1233] = !f[633] && f[683] && !f[156]; // c0t860i86
	assign leaf[1234] = !f[633] && f[683] && f[156] && !f[235]; // c0t860i86
	assign leaf[1235] = !f[633] && f[683] && f[156] && f[235]; // c0t860i86
	assign leaf[1236] = f[633] && !f[579] && !f[576]; // c0t860i86
	assign leaf[1237] = f[633] && !f[579] && f[576] && !f[542]; // c0t860i86
	assign leaf[1238] = f[633] && !f[579] && f[576] && f[542]; // c0t860i86
	assign leaf[1239] = f[633] && f[579] && !f[234] && !f[266]; // c0t860i86
	assign leaf[1240] = f[633] && f[579] && !f[234] && f[266]; // c0t860i86
	assign leaf[1241] = f[633] && f[579] && f[234] && !f[157]; // c0t860i86
	assign leaf[1242] = f[633] && f[579] && f[234] && f[157]; // c0t860i86
	assign leaf[1243] = !f[380] && !f[456] && !f[516] && !f[212]; // c0t870i87
	assign leaf[1244] = !f[380] && !f[456] && !f[516] && f[212]; // c0t870i87
	assign leaf[1245] = !f[380] && !f[456] && f[516] && !f[266]; // c0t870i87
	assign leaf[1246] = !f[380] && !f[456] && f[516] && f[266]; // c0t870i87
	assign leaf[1247] = !f[380] && f[456] && !f[654] && !f[520]; // c0t870i87
	assign leaf[1248] = !f[380] && f[456] && !f[654] && f[520]; // c0t870i87
	assign leaf[1249] = !f[380] && f[456] && f[654] && !f[681]; // c0t870i87
	assign leaf[1250] = !f[380] && f[456] && f[654] && f[681]; // c0t870i87
	assign leaf[1251] = f[380] && !f[378] && !f[377] && !f[412]; // c0t870i87
	assign leaf[1252] = f[380] && !f[378] && !f[377] && f[412]; // c0t870i87
	assign leaf[1253] = f[380] && !f[378] && f[377]; // c0t870i87
	assign leaf[1254] = f[380] && f[378] && !f[427] && !f[410]; // c0t870i87
	assign leaf[1255] = f[380] && f[378] && !f[427] && f[410]; // c0t870i87
	assign leaf[1256] = f[380] && f[378] && f[427] && !f[273]; // c0t870i87
	assign leaf[1257] = f[380] && f[378] && f[427] && f[273]; // c0t870i87
	assign leaf[1258] = !f[514] && !f[539] && !f[513] && !f[508]; // c0t880i88
	assign leaf[1259] = !f[514] && !f[539] && !f[513] && f[508]; // c0t880i88
	assign leaf[1260] = !f[514] && !f[539] && f[513] && !f[185]; // c0t880i88
	assign leaf[1261] = !f[514] && !f[539] && f[513] && f[185]; // c0t880i88
	assign leaf[1262] = !f[514] && f[539] && !f[624] && !f[183]; // c0t880i88
	assign leaf[1263] = !f[514] && f[539] && !f[624] && f[183]; // c0t880i88
	assign leaf[1264] = !f[514] && f[539] && f[624] && !f[483]; // c0t880i88
	assign leaf[1265] = !f[514] && f[539] && f[624] && f[483]; // c0t880i88
	assign leaf[1266] = f[514] && !f[567] && !f[465] && !f[349]; // c0t880i88
	assign leaf[1267] = f[514] && !f[567] && !f[465] && f[349]; // c0t880i88
	assign leaf[1268] = f[514] && !f[567] && f[465] && !f[268]; // c0t880i88
	assign leaf[1269] = f[514] && !f[567] && f[465] && f[268]; // c0t880i88
	assign leaf[1270] = f[514] && f[567] && !f[371] && !f[651]; // c0t880i88
	assign leaf[1271] = f[514] && f[567] && !f[371] && f[651]; // c0t880i88
	assign leaf[1272] = f[514] && f[567] && f[371]; // c0t880i88
	assign leaf[1273] = !f[602] && !f[456] && !f[687] && !f[356]; // c0t890i89
	assign leaf[1274] = !f[602] && !f[456] && !f[687] && f[356]; // c0t890i89
	assign leaf[1275] = !f[602] && !f[456] && f[687] && !f[156]; // c0t890i89
	assign leaf[1276] = !f[602] && !f[456] && f[687] && f[156]; // c0t890i89
	assign leaf[1277] = !f[602] && f[456] && !f[356] && !f[598]; // c0t890i89
	assign leaf[1278] = !f[602] && f[456] && !f[356] && f[598]; // c0t890i89
	assign leaf[1279] = !f[602] && f[456] && f[356] && !f[433]; // c0t890i89
	assign leaf[1280] = !f[602] && f[456] && f[356] && f[433]; // c0t890i89
	assign leaf[1281] = f[602] && !f[128] && !f[491] && !f[372]; // c0t890i89
	assign leaf[1282] = f[602] && !f[128] && !f[491] && f[372]; // c0t890i89
	assign leaf[1283] = f[602] && !f[128] && f[491] && !f[596]; // c0t890i89
	assign leaf[1284] = f[602] && !f[128] && f[491] && f[596]; // c0t890i89
	assign leaf[1285] = f[602] && f[128] && !f[322] && !f[435]; // c0t890i89
	assign leaf[1286] = f[602] && f[128] && !f[322] && f[435]; // c0t890i89
	assign leaf[1287] = f[602] && f[128] && f[322] && !f[463]; // c0t890i89
	assign leaf[1288] = f[602] && f[128] && f[322] && f[463]; // c0t890i89
	assign leaf[1289] = !f[240] && !f[325] && !f[214] && !f[331]; // c0t900i90
	assign leaf[1290] = !f[240] && !f[325] && !f[214] && f[331]; // c0t900i90
	assign leaf[1291] = !f[240] && !f[325] && f[214] && !f[128]; // c0t900i90
	assign leaf[1292] = !f[240] && !f[325] && f[214] && f[128]; // c0t900i90
	assign leaf[1293] = !f[240] && f[325] && !f[460] && !f[370]; // c0t900i90
	assign leaf[1294] = !f[240] && f[325] && !f[460] && f[370]; // c0t900i90
	assign leaf[1295] = !f[240] && f[325] && f[460]; // c0t900i90
	assign leaf[1296] = f[240] && !f[466] && !f[374] && !f[511]; // c0t900i90
	assign leaf[1297] = f[240] && !f[466] && !f[374] && f[511]; // c0t900i90
	assign leaf[1298] = f[240] && !f[466] && f[374] && !f[468]; // c0t900i90
	assign leaf[1299] = f[240] && !f[466] && f[374] && f[468]; // c0t900i90
	assign leaf[1300] = f[240] && f[466] && !f[403] && !f[400]; // c0t900i90
	assign leaf[1301] = f[240] && f[466] && !f[403] && f[400]; // c0t900i90
	assign leaf[1302] = f[240] && f[466] && f[403] && !f[457]; // c0t900i90
	assign leaf[1303] = f[240] && f[466] && f[403] && f[457]; // c0t900i90
	assign leaf[1304] = !f[663] && !f[583] && !f[513] && !f[328]; // c0t910i91
	assign leaf[1305] = !f[663] && !f[583] && !f[513] && f[328]; // c0t910i91
	assign leaf[1306] = !f[663] && !f[583] && f[513] && !f[183]; // c0t910i91
	assign leaf[1307] = !f[663] && !f[583] && f[513] && f[183]; // c0t910i91
	assign leaf[1308] = !f[663] && f[583]; // c0t910i91
	assign leaf[1309] = f[663] && !f[346]; // c0t910i91
	assign leaf[1310] = f[663] && f[346]; // c0t910i91
	assign leaf[1311] = !f[605] && !f[260] && !f[242] && !f[566]; // c0t920i92
	assign leaf[1312] = !f[605] && !f[260] && !f[242] && f[566]; // c0t920i92
	assign leaf[1313] = !f[605] && !f[260] && f[242] && !f[683]; // c0t920i92
	assign leaf[1314] = !f[605] && !f[260] && f[242] && f[683]; // c0t920i92
	assign leaf[1315] = !f[605] && f[260] && !f[359] && !f[545]; // c0t920i92
	assign leaf[1316] = !f[605] && f[260] && !f[359] && f[545]; // c0t920i92
	assign leaf[1317] = !f[605] && f[260] && f[359]; // c0t920i92
	assign leaf[1318] = f[605] && !f[397] && !f[597] && !f[599]; // c0t920i92
	assign leaf[1319] = f[605] && !f[397] && !f[597] && f[599]; // c0t920i92
	assign leaf[1320] = f[605] && !f[397] && f[597] && !f[484]; // c0t920i92
	assign leaf[1321] = f[605] && !f[397] && f[597] && f[484]; // c0t920i92
	assign leaf[1322] = f[605] && f[397] && !f[207]; // c0t920i92
	assign leaf[1323] = f[605] && f[397] && f[207] && !f[428]; // c0t920i92
	assign leaf[1324] = f[605] && f[397] && f[207] && f[428]; // c0t920i92
	assign leaf[1325] = !f[294] && !f[351] && !f[518] && !f[344]; // c0t930i93
	assign leaf[1326] = !f[294] && !f[351] && !f[518] && f[344]; // c0t930i93
	assign leaf[1327] = !f[294] && !f[351] && f[518] && !f[455]; // c0t930i93
	assign leaf[1328] = !f[294] && !f[351] && f[518] && f[455]; // c0t930i93
	assign leaf[1329] = !f[294] && f[351] && !f[376]; // c0t930i93
	assign leaf[1330] = !f[294] && f[351] && f[376]; // c0t930i93
	assign leaf[1331] = f[294] && !f[99] && !f[384] && !f[160]; // c0t930i93
	assign leaf[1332] = f[294] && !f[99] && !f[384] && f[160]; // c0t930i93
	assign leaf[1333] = f[294] && !f[99] && f[384] && !f[402]; // c0t930i93
	assign leaf[1334] = f[294] && !f[99] && f[384] && f[402]; // c0t930i93
	assign leaf[1335] = f[294] && f[99]; // c0t930i93
	assign leaf[1336] = !f[434] && !f[526] && !f[319] && !f[291]; // c0t940i94
	assign leaf[1337] = !f[434] && !f[526] && !f[319] && f[291]; // c0t940i94
	assign leaf[1338] = !f[434] && !f[526] && f[319] && !f[468]; // c0t940i94
	assign leaf[1339] = !f[434] && !f[526] && f[319] && f[468]; // c0t940i94
	assign leaf[1340] = !f[434] && f[526] && !f[427] && !f[413]; // c0t940i94
	assign leaf[1341] = !f[434] && f[526] && !f[427] && f[413]; // c0t940i94
	assign leaf[1342] = !f[434] && f[526] && f[427] && !f[208]; // c0t940i94
	assign leaf[1343] = !f[434] && f[526] && f[427] && f[208]; // c0t940i94
	assign leaf[1344] = f[434] && !f[273] && !f[316]; // c0t940i94
	assign leaf[1345] = f[434] && !f[273] && f[316]; // c0t940i94
	assign leaf[1346] = f[434] && f[273] && !f[349]; // c0t940i94
	assign leaf[1347] = f[434] && f[273] && f[349] && !f[595]; // c0t940i94
	assign leaf[1348] = f[434] && f[273] && f[349] && f[595]; // c0t940i94
	assign leaf[1349] = !f[408] && !f[574] && !f[233] && !f[541]; // c0t950i95
	assign leaf[1350] = !f[408] && !f[574] && !f[233] && f[541]; // c0t950i95
	assign leaf[1351] = !f[408] && !f[574] && f[233] && !f[347]; // c0t950i95
	assign leaf[1352] = !f[408] && !f[574] && f[233] && f[347]; // c0t950i95
	assign leaf[1353] = !f[408] && f[574] && !f[354] && !f[190]; // c0t950i95
	assign leaf[1354] = !f[408] && f[574] && !f[354] && f[190]; // c0t950i95
	assign leaf[1355] = !f[408] && f[574] && f[354] && !f[240]; // c0t950i95
	assign leaf[1356] = !f[408] && f[574] && f[354] && f[240]; // c0t950i95
	assign leaf[1357] = f[408] && !f[464] && !f[600]; // c0t950i95
	assign leaf[1358] = f[408] && !f[464] && f[600]; // c0t950i95
	assign leaf[1359] = f[408] && f[464] && !f[571]; // c0t950i95
	assign leaf[1360] = f[408] && f[464] && f[571] && !f[577]; // c0t950i95
	assign leaf[1361] = f[408] && f[464] && f[571] && f[577]; // c0t950i95
	assign leaf[1362] = !f[294] && !f[547] && !f[659] && !f[550]; // c0t960i96
	assign leaf[1363] = !f[294] && !f[547] && !f[659] && f[550]; // c0t960i96
	assign leaf[1364] = !f[294] && !f[547] && f[659] && !f[432]; // c0t960i96
	assign leaf[1365] = !f[294] && !f[547] && f[659] && f[432]; // c0t960i96
	assign leaf[1366] = !f[294] && f[547] && !f[660] && !f[599]; // c0t960i96
	assign leaf[1367] = !f[294] && f[547] && !f[660] && f[599]; // c0t960i96
	assign leaf[1368] = !f[294] && f[547] && f[660]; // c0t960i96
	assign leaf[1369] = f[294] && !f[435] && !f[331] && !f[327]; // c0t960i96
	assign leaf[1370] = f[294] && !f[435] && !f[331] && f[327]; // c0t960i96
	assign leaf[1371] = f[294] && !f[435] && f[331] && !f[539]; // c0t960i96
	assign leaf[1372] = f[294] && !f[435] && f[331] && f[539]; // c0t960i96
	assign leaf[1373] = f[294] && f[435] && !f[434] && !f[244]; // c0t960i96
	assign leaf[1374] = f[294] && f[435] && !f[434] && f[244]; // c0t960i96
	assign leaf[1375] = f[294] && f[435] && f[434] && !f[130]; // c0t960i96
	assign leaf[1376] = f[294] && f[435] && f[434] && f[130]; // c0t960i96
	assign leaf[1377] = !f[555] && !f[468] && !f[602] && !f[460]; // c0t970i97
	assign leaf[1378] = !f[555] && !f[468] && !f[602] && f[460]; // c0t970i97
	assign leaf[1379] = !f[555] && !f[468] && f[602] && !f[432]; // c0t970i97
	assign leaf[1380] = !f[555] && !f[468] && f[602] && f[432]; // c0t970i97
	assign leaf[1381] = !f[555] && f[468] && !f[295] && !f[268]; // c0t970i97
	assign leaf[1382] = !f[555] && f[468] && !f[295] && f[268]; // c0t970i97
	assign leaf[1383] = !f[555] && f[468] && f[295] && !f[569]; // c0t970i97
	assign leaf[1384] = !f[555] && f[468] && f[295] && f[569]; // c0t970i97
	assign leaf[1385] = f[555] && !f[398]; // c0t970i97
	assign leaf[1386] = f[555] && f[398]; // c0t970i97
	assign leaf[1387] = !f[425] && !f[542] && !f[541] && !f[271]; // c0t980i98
	assign leaf[1388] = !f[425] && !f[542] && !f[541] && f[271]; // c0t980i98
	assign leaf[1389] = !f[425] && !f[542] && f[541] && !f[382]; // c0t980i98
	assign leaf[1390] = !f[425] && !f[542] && f[541] && f[382]; // c0t980i98
	assign leaf[1391] = !f[425] && f[542] && !f[247] && !f[510]; // c0t980i98
	assign leaf[1392] = !f[425] && f[542] && !f[247] && f[510]; // c0t980i98
	assign leaf[1393] = !f[425] && f[542] && f[247]; // c0t980i98
	assign leaf[1394] = f[425] && !f[471] && !f[396] && !f[343]; // c0t980i98
	assign leaf[1395] = f[425] && !f[471] && !f[396] && f[343]; // c0t980i98
	assign leaf[1396] = f[425] && !f[471] && f[396]; // c0t980i98
	assign leaf[1397] = f[425] && f[471] && !f[317]; // c0t980i98
	assign leaf[1398] = f[425] && f[471] && f[317]; // c0t980i98
	assign leaf[1399] = !f[386] && !f[354] && !f[416] && !f[356]; // c0t990i99
	assign leaf[1400] = !f[386] && !f[354] && !f[416] && f[356]; // c0t990i99
	assign leaf[1401] = !f[386] && !f[354] && f[416]; // c0t990i99
	assign leaf[1402] = !f[386] && f[354] && !f[187] && !f[515]; // c0t990i99
	assign leaf[1403] = !f[386] && f[354] && !f[187] && f[515]; // c0t990i99
	assign leaf[1404] = !f[386] && f[354] && f[187] && !f[130]; // c0t990i99
	assign leaf[1405] = !f[386] && f[354] && f[187] && f[130]; // c0t990i99
	assign leaf[1406] = f[386] && !f[159] && !f[383] && !f[273]; // c0t990i99
	assign leaf[1407] = f[386] && !f[159] && !f[383] && f[273]; // c0t990i99
	assign leaf[1408] = f[386] && !f[159] && f[383] && !f[297]; // c0t990i99
	assign leaf[1409] = f[386] && !f[159] && f[383] && f[297]; // c0t990i99
	assign leaf[1410] = f[386] && f[159] && !f[570]; // c0t990i99
	assign leaf[1411] = f[386] && f[159] && f[570]; // c0t990i99
endmodule

module decision_tree_leaves_1(input logic [0:783] f, output logic [0:1154] leaf);
	assign leaf[0] = !f[350] && !f[351] && !f[349]; // c1t1i0
	assign leaf[1] = !f[350] && !f[351] && f[349] && !f[347]; // c1t1i0
	assign leaf[2] = !f[350] && !f[351] && f[349] && f[347]; // c1t1i0
	assign leaf[3] = !f[350] && f[351] && !f[236] && !f[492]; // c1t1i0
	assign leaf[4] = !f[350] && f[351] && !f[236] && f[492]; // c1t1i0
	assign leaf[5] = !f[350] && f[351] && f[236] && !f[608]; // c1t1i0
	assign leaf[6] = !f[350] && f[351] && f[236] && f[608]; // c1t1i0
	assign leaf[7] = f[350] && !f[489] && !f[490] && !f[488]; // c1t1i0
	assign leaf[8] = f[350] && !f[489] && !f[490] && f[488]; // c1t1i0
	assign leaf[9] = f[350] && !f[489] && f[490] && !f[404]; // c1t1i0
	assign leaf[10] = f[350] && !f[489] && f[490] && f[404]; // c1t1i0
	assign leaf[11] = f[350] && f[489] && !f[521] && !f[375]; // c1t1i0
	assign leaf[12] = f[350] && f[489] && !f[521] && f[375]; // c1t1i0
	assign leaf[13] = f[350] && f[489] && f[521] && !f[487]; // c1t1i0
	assign leaf[14] = f[350] && f[489] && f[521] && f[487]; // c1t1i0
	assign leaf[15] = !f[409] && !f[378] && !f[379] && !f[377]; // c1t11i1
	assign leaf[16] = !f[409] && !f[378] && !f[379] && f[377]; // c1t11i1
	assign leaf[17] = !f[409] && !f[378] && f[379] && !f[353]; // c1t11i1
	assign leaf[18] = !f[409] && !f[378] && f[379] && f[353]; // c1t11i1
	assign leaf[19] = !f[409] && f[378] && !f[550] && !f[319]; // c1t11i1
	assign leaf[20] = !f[409] && f[378] && !f[550] && f[319]; // c1t11i1
	assign leaf[21] = !f[409] && f[378] && f[550] && !f[293]; // c1t11i1
	assign leaf[22] = !f[409] && f[378] && f[550] && f[293]; // c1t11i1
	assign leaf[23] = f[409] && !f[410] && !f[323] && !f[594]; // c1t11i1
	assign leaf[24] = f[409] && !f[410] && !f[323] && f[594]; // c1t11i1
	assign leaf[25] = f[409] && !f[410] && f[323] && !f[544]; // c1t11i1
	assign leaf[26] = f[409] && !f[410] && f[323] && f[544]; // c1t11i1
	assign leaf[27] = f[409] && f[410] && !f[171] && !f[613]; // c1t11i1
	assign leaf[28] = f[409] && f[410] && !f[171] && f[613]; // c1t11i1
	assign leaf[29] = f[409] && f[410] && f[171]; // c1t11i1
	assign leaf[30] = !f[437] && !f[262] && !f[406] && !f[407]; // c1t21i2
	assign leaf[31] = !f[437] && !f[262] && !f[406] && f[407]; // c1t21i2
	assign leaf[32] = !f[437] && !f[262] && f[406] && !f[178]; // c1t21i2
	assign leaf[33] = !f[437] && !f[262] && f[406] && f[178]; // c1t21i2
	assign leaf[34] = !f[437] && f[262] && !f[325] && !f[350]; // c1t21i2
	assign leaf[35] = !f[437] && f[262] && !f[325] && f[350]; // c1t21i2
	assign leaf[36] = !f[437] && f[262] && f[325]; // c1t21i2
	assign leaf[37] = f[437] && !f[438] && !f[322] && !f[622]; // c1t21i2
	assign leaf[38] = f[437] && !f[438] && !f[322] && f[622]; // c1t21i2
	assign leaf[39] = f[437] && !f[438] && f[322] && !f[545]; // c1t21i2
	assign leaf[40] = f[437] && !f[438] && f[322] && f[545]; // c1t21i2
	assign leaf[41] = f[437] && f[438] && !f[613] && !f[69]; // c1t21i2
	assign leaf[42] = f[437] && f[438] && !f[613] && f[69]; // c1t21i2
	assign leaf[43] = f[437] && f[438] && f[613]; // c1t21i2
	assign leaf[44] = !f[350] && !f[351] && !f[382] && !f[374]; // c1t31i3
	assign leaf[45] = !f[350] && !f[351] && !f[382] && f[374]; // c1t31i3
	assign leaf[46] = !f[350] && !f[351] && f[382]; // c1t31i3
	assign leaf[47] = !f[350] && f[351] && !f[209] && !f[431]; // c1t31i3
	assign leaf[48] = !f[350] && f[351] && !f[209] && f[431]; // c1t31i3
	assign leaf[49] = !f[350] && f[351] && f[209] && !f[406]; // c1t31i3
	assign leaf[50] = !f[350] && f[351] && f[209] && f[406]; // c1t31i3
	assign leaf[51] = f[350] && !f[375] && !f[234] && !f[327]; // c1t31i3
	assign leaf[52] = f[350] && !f[375] && !f[234] && f[327]; // c1t31i3
	assign leaf[53] = f[350] && !f[375] && f[234] && !f[297]; // c1t31i3
	assign leaf[54] = f[350] && !f[375] && f[234] && f[297]; // c1t31i3
	assign leaf[55] = f[350] && f[375] && !f[374] && !f[517]; // c1t31i3
	assign leaf[56] = f[350] && f[375] && !f[374] && f[517]; // c1t31i3
	assign leaf[57] = f[350] && f[375] && f[374] && !f[294]; // c1t31i3
	assign leaf[58] = f[350] && f[375] && f[374] && f[294]; // c1t31i3
	assign leaf[59] = !f[437] && !f[346] && !f[578] && !f[300]; // c1t41i4
	assign leaf[60] = !f[437] && !f[346] && !f[578] && f[300]; // c1t41i4
	assign leaf[61] = !f[437] && !f[346] && f[578] && !f[293]; // c1t41i4
	assign leaf[62] = !f[437] && !f[346] && f[578] && f[293]; // c1t41i4
	assign leaf[63] = !f[437] && f[346] && !f[294] && !f[120]; // c1t41i4
	assign leaf[64] = !f[437] && f[346] && !f[294] && f[120]; // c1t41i4
	assign leaf[65] = !f[437] && f[346] && f[294] && !f[435]; // c1t41i4
	assign leaf[66] = !f[437] && f[346] && f[294] && f[435]; // c1t41i4
	assign leaf[67] = f[437] && !f[438] && !f[323] && !f[436]; // c1t41i4
	assign leaf[68] = f[437] && !f[438] && !f[323] && f[436]; // c1t41i4
	assign leaf[69] = f[437] && !f[438] && f[323] && !f[489]; // c1t41i4
	assign leaf[70] = f[437] && !f[438] && f[323] && f[489]; // c1t41i4
	assign leaf[71] = f[437] && f[438] && !f[69]; // c1t41i4
	assign leaf[72] = f[437] && f[438] && f[69] && !f[383]; // c1t41i4
	assign leaf[73] = f[437] && f[438] && f[69] && f[383]; // c1t41i4
	assign leaf[74] = !f[382] && !f[465] && !f[378] && !f[379]; // c1t51i5
	assign leaf[75] = !f[382] && !f[465] && !f[378] && f[379]; // c1t51i5
	assign leaf[76] = !f[382] && !f[465] && f[378] && !f[206]; // c1t51i5
	assign leaf[77] = !f[382] && !f[465] && f[378] && f[206]; // c1t51i5
	assign leaf[78] = !f[382] && f[465] && !f[466] && !f[518]; // c1t51i5
	assign leaf[79] = !f[382] && f[465] && !f[466] && f[518]; // c1t51i5
	assign leaf[80] = !f[382] && f[465] && f[466] && !f[98]; // c1t51i5
	assign leaf[81] = !f[382] && f[465] && f[466] && f[98]; // c1t51i5
	assign leaf[82] = f[382] && !f[162] && !f[355] && !f[488]; // c1t51i5
	assign leaf[83] = f[382] && !f[162] && !f[355] && f[488]; // c1t51i5
	assign leaf[84] = f[382] && !f[162] && f[355]; // c1t51i5
	assign leaf[85] = f[382] && f[162] && !f[269] && !f[296]; // c1t51i5
	assign leaf[86] = f[382] && f[162] && !f[269] && f[296]; // c1t51i5
	assign leaf[87] = f[382] && f[162] && f[269] && !f[320]; // c1t51i5
	assign leaf[88] = f[382] && f[162] && f[269] && f[320]; // c1t51i5
	assign leaf[89] = !f[323] && !f[322] && !f[211] && !f[650]; // c1t61i6
	assign leaf[90] = !f[323] && !f[322] && !f[211] && f[650]; // c1t61i6
	assign leaf[91] = !f[323] && !f[322] && f[211] && !f[378]; // c1t61i6
	assign leaf[92] = !f[323] && !f[322] && f[211] && f[378]; // c1t61i6
	assign leaf[93] = !f[323] && f[322] && !f[627] && !f[380]; // c1t61i6
	assign leaf[94] = !f[323] && f[322] && !f[627] && f[380]; // c1t61i6
	assign leaf[95] = !f[323] && f[322] && f[627] && !f[126]; // c1t61i6
	assign leaf[96] = !f[323] && f[322] && f[627] && f[126]; // c1t61i6
	assign leaf[97] = f[323] && !f[494] && !f[234] && !f[402]; // c1t61i6
	assign leaf[98] = f[323] && !f[494] && !f[234] && f[402]; // c1t61i6
	assign leaf[99] = f[323] && !f[494] && f[234] && !f[324]; // c1t61i6
	assign leaf[100] = f[323] && !f[494] && f[234] && f[324]; // c1t61i6
	assign leaf[101] = f[323] && f[494] && !f[71] && !f[98]; // c1t61i6
	assign leaf[102] = f[323] && f[494] && !f[71] && f[98]; // c1t61i6
	assign leaf[103] = f[323] && f[494] && f[71]; // c1t61i6
	assign leaf[104] = !f[323] && !f[212] && !f[322] && !f[650]; // c1t71i7
	assign leaf[105] = !f[323] && !f[212] && !f[322] && f[650]; // c1t71i7
	assign leaf[106] = !f[323] && !f[212] && f[322] && !f[380]; // c1t71i7
	assign leaf[107] = !f[323] && !f[212] && f[322] && f[380]; // c1t71i7
	assign leaf[108] = !f[323] && f[212] && !f[406] && !f[620]; // c1t71i7
	assign leaf[109] = !f[323] && f[212] && !f[406] && f[620]; // c1t71i7
	assign leaf[110] = !f[323] && f[212] && f[406] && !f[437]; // c1t71i7
	assign leaf[111] = !f[323] && f[212] && f[406] && f[437]; // c1t71i7
	assign leaf[112] = f[323] && !f[430] && !f[434] && !f[349]; // c1t71i7
	assign leaf[113] = f[323] && !f[430] && !f[434] && f[349]; // c1t71i7
	assign leaf[114] = f[323] && !f[430] && f[434] && !f[205]; // c1t71i7
	assign leaf[115] = f[323] && !f[430] && f[434] && f[205]; // c1t71i7
	assign leaf[116] = f[323] && f[430] && !f[236] && !f[189]; // c1t71i7
	assign leaf[117] = f[323] && f[430] && !f[236] && f[189]; // c1t71i7
	assign leaf[118] = f[323] && f[430] && f[236] && !f[347]; // c1t71i7
	assign leaf[119] = f[323] && f[430] && f[236] && f[347]; // c1t71i7
	assign leaf[120] = !f[402] && !f[406] && !f[99] && !f[405]; // c1t81i8
	assign leaf[121] = !f[402] && !f[406] && !f[99] && f[405]; // c1t81i8
	assign leaf[122] = !f[402] && !f[406] && f[99] && !f[379]; // c1t81i8
	assign leaf[123] = !f[402] && !f[406] && f[99] && f[379]; // c1t81i8
	assign leaf[124] = !f[402] && f[406] && !f[233] && !f[295]; // c1t81i8
	assign leaf[125] = !f[402] && f[406] && !f[233] && f[295]; // c1t81i8
	assign leaf[126] = !f[402] && f[406] && f[233] && !f[269]; // c1t81i8
	assign leaf[127] = !f[402] && f[406] && f[233] && f[269]; // c1t81i8
	assign leaf[128] = f[402] && !f[295]; // c1t81i8
	assign leaf[129] = f[402] && f[295] && !f[494] && !f[373]; // c1t81i8
	assign leaf[130] = f[402] && f[295] && !f[494] && f[373]; // c1t81i8
	assign leaf[131] = f[402] && f[295] && f[494]; // c1t81i8
	assign leaf[132] = !f[410] && !f[318] && !f[511] && !f[205]; // c1t91i9
	assign leaf[133] = !f[410] && !f[318] && !f[511] && f[205]; // c1t91i9
	assign leaf[134] = !f[410] && !f[318] && f[511] && !f[649]; // c1t91i9
	assign leaf[135] = !f[410] && !f[318] && f[511] && f[649]; // c1t91i9
	assign leaf[136] = !f[410] && f[318] && !f[294] && !f[148]; // c1t91i9
	assign leaf[137] = !f[410] && f[318] && !f[294] && f[148]; // c1t91i9
	assign leaf[138] = !f[410] && f[318] && f[294] && !f[126]; // c1t91i9
	assign leaf[139] = !f[410] && f[318] && f[294] && f[126]; // c1t91i9
	assign leaf[140] = f[410] && !f[163] && !f[411] && !f[322]; // c1t91i9
	assign leaf[141] = f[410] && !f[163] && !f[411] && f[322]; // c1t91i9
	assign leaf[142] = f[410] && !f[163] && f[411]; // c1t91i9
	assign leaf[143] = f[410] && f[163] && !f[269]; // c1t91i9
	assign leaf[144] = f[410] && f[163] && f[269]; // c1t91i9
	assign leaf[145] = !f[430] && !f[434] && !f[433] && !f[101]; // c1t101i10
	assign leaf[146] = !f[430] && !f[434] && !f[433] && f[101]; // c1t101i10
	assign leaf[147] = !f[430] && !f[434] && f[433] && !f[548]; // c1t101i10
	assign leaf[148] = !f[430] && !f[434] && f[433] && f[548]; // c1t101i10
	assign leaf[149] = !f[430] && f[434] && !f[299] && !f[322]; // c1t101i10
	assign leaf[150] = !f[430] && f[434] && !f[299] && f[322]; // c1t101i10
	assign leaf[151] = !f[430] && f[434] && f[299] && !f[183]; // c1t101i10
	assign leaf[152] = !f[430] && f[434] && f[299] && f[183]; // c1t101i10
	assign leaf[153] = f[430] && !f[349] && !f[649] && !f[743]; // c1t101i10
	assign leaf[154] = f[430] && !f[349] && !f[649] && f[743]; // c1t101i10
	assign leaf[155] = f[430] && !f[349] && f[649] && !f[184]; // c1t101i10
	assign leaf[156] = f[430] && !f[349] && f[649] && f[184]; // c1t101i10
	assign leaf[157] = f[430] && f[349] && !f[521] && !f[268]; // c1t101i10
	assign leaf[158] = f[430] && f[349] && !f[521] && f[268]; // c1t101i10
	assign leaf[159] = f[430] && f[349] && f[521]; // c1t101i10
	assign leaf[160] = !f[466] && !f[374] && !f[511] && !f[683]; // c1t111i11
	assign leaf[161] = !f[466] && !f[374] && !f[511] && f[683]; // c1t111i11
	assign leaf[162] = !f[466] && !f[374] && f[511] && !f[649]; // c1t111i11
	assign leaf[163] = !f[466] && !f[374] && f[511] && f[649]; // c1t111i11
	assign leaf[164] = !f[466] && f[374] && !f[294]; // c1t111i11
	assign leaf[165] = !f[466] && f[374] && f[294] && !f[404]; // c1t111i11
	assign leaf[166] = !f[466] && f[374] && f[294] && f[404]; // c1t111i11
	assign leaf[167] = f[466] && !f[145] && !f[556] && !f[467]; // c1t111i11
	assign leaf[168] = f[466] && !f[145] && !f[556] && f[467]; // c1t111i11
	assign leaf[169] = f[466] && !f[145] && f[556]; // c1t111i11
	assign leaf[170] = f[466] && f[145]; // c1t111i11
	assign leaf[171] = !f[438] && !f[235] && !f[493] && !f[150]; // c1t121i12
	assign leaf[172] = !f[438] && !f[235] && !f[493] && f[150]; // c1t121i12
	assign leaf[173] = !f[438] && !f[235] && f[493] && !f[181]; // c1t121i12
	assign leaf[174] = !f[438] && !f[235] && f[493] && f[181]; // c1t121i12
	assign leaf[175] = !f[438] && f[235] && !f[151] && !f[98]; // c1t121i12
	assign leaf[176] = !f[438] && f[235] && !f[151] && f[98]; // c1t121i12
	assign leaf[177] = !f[438] && f[235] && f[151] && !f[265]; // c1t121i12
	assign leaf[178] = !f[438] && f[235] && f[151] && f[265]; // c1t121i12
	assign leaf[179] = f[438] && !f[439] && !f[609] && !f[123]; // c1t121i12
	assign leaf[180] = f[438] && !f[439] && !f[609] && f[123]; // c1t121i12
	assign leaf[181] = f[438] && !f[439] && f[609]; // c1t121i12
	assign leaf[182] = f[438] && f[439] && !f[163]; // c1t121i12
	assign leaf[183] = f[438] && f[439] && f[163]; // c1t121i12
	assign leaf[184] = !f[429] && !f[354] && !f[272] && !f[462]; // c1t131i13
	assign leaf[185] = !f[429] && !f[354] && !f[272] && f[462]; // c1t131i13
	assign leaf[186] = !f[429] && !f[354] && f[272] && !f[518]; // c1t131i13
	assign leaf[187] = !f[429] && !f[354] && f[272] && f[518]; // c1t131i13
	assign leaf[188] = !f[429] && f[354] && !f[162] && !f[296]; // c1t131i13
	assign leaf[189] = !f[429] && f[354] && !f[162] && f[296]; // c1t131i13
	assign leaf[190] = !f[429] && f[354] && f[162] && !f[211]; // c1t131i13
	assign leaf[191] = !f[429] && f[354] && f[162] && f[211]; // c1t131i13
	assign leaf[192] = f[429] && !f[375]; // c1t131i13
	assign leaf[193] = f[429] && f[375] && !f[687] && !f[679]; // c1t131i13
	assign leaf[194] = f[429] && f[375] && !f[687] && f[679]; // c1t131i13
	assign leaf[195] = f[429] && f[375] && f[687] && !f[345]; // c1t131i13
	assign leaf[196] = f[429] && f[375] && f[687] && f[345]; // c1t131i13
	assign leaf[197] = !f[355] && !f[684] && !f[467] && !f[510]; // c1t141i14
	assign leaf[198] = !f[355] && !f[684] && !f[467] && f[510]; // c1t141i14
	assign leaf[199] = !f[355] && !f[684] && f[467] && !f[98]; // c1t141i14
	assign leaf[200] = !f[355] && !f[684] && f[467] && f[98]; // c1t141i14
	assign leaf[201] = !f[355] && f[684] && !f[208] && !f[295]; // c1t141i14
	assign leaf[202] = !f[355] && f[684] && !f[208] && f[295]; // c1t141i14
	assign leaf[203] = !f[355] && f[684] && f[208] && !f[409]; // c1t141i14
	assign leaf[204] = !f[355] && f[684] && f[208] && f[409]; // c1t141i14
	assign leaf[205] = f[355] && !f[161] && !f[192] && !f[102]; // c1t141i14
	assign leaf[206] = f[355] && !f[161] && !f[192] && f[102]; // c1t141i14
	assign leaf[207] = f[355] && !f[161] && f[192]; // c1t141i14
	assign leaf[208] = f[355] && f[161] && !f[211] && !f[651]; // c1t141i14
	assign leaf[209] = f[355] && f[161] && !f[211] && f[651]; // c1t141i14
	assign leaf[210] = f[355] && f[161] && f[211] && !f[659]; // c1t141i14
	assign leaf[211] = f[355] && f[161] && f[211] && f[659]; // c1t141i14
	assign leaf[212] = !f[430] && !f[434] && !f[100] && !f[189]; // c1t151i15
	assign leaf[213] = !f[430] && !f[434] && !f[100] && f[189]; // c1t151i15
	assign leaf[214] = !f[430] && !f[434] && f[100] && !f[350]; // c1t151i15
	assign leaf[215] = !f[430] && !f[434] && f[100] && f[350]; // c1t151i15
	assign leaf[216] = !f[430] && f[434] && !f[298] && !f[486]; // c1t151i15
	assign leaf[217] = !f[430] && f[434] && !f[298] && f[486]; // c1t151i15
	assign leaf[218] = !f[430] && f[434] && f[298] && !f[237]; // c1t151i15
	assign leaf[219] = !f[430] && f[434] && f[298] && f[237]; // c1t151i15
	assign leaf[220] = f[430] && !f[349] && !f[649] && !f[715]; // c1t151i15
	assign leaf[221] = f[430] && !f[349] && !f[649] && f[715]; // c1t151i15
	assign leaf[222] = f[430] && !f[349] && f[649]; // c1t151i15
	assign leaf[223] = f[430] && f[349] && !f[408] && !f[519]; // c1t151i15
	assign leaf[224] = f[430] && f[349] && !f[408] && f[519]; // c1t151i15
	assign leaf[225] = f[430] && f[349] && f[408] && !f[410]; // c1t151i15
	assign leaf[226] = f[430] && f[349] && f[408] && f[410]; // c1t151i15
	assign leaf[227] = !f[317] && !f[628] && !f[684] && !f[204]; // c1t161i16
	assign leaf[228] = !f[317] && !f[628] && !f[684] && f[204]; // c1t161i16
	assign leaf[229] = !f[317] && !f[628] && f[684] && !f[631]; // c1t161i16
	assign leaf[230] = !f[317] && !f[628] && f[684] && f[631]; // c1t161i16
	assign leaf[231] = !f[317] && f[628] && !f[545] && !f[405]; // c1t161i16
	assign leaf[232] = !f[317] && f[628] && !f[545] && f[405]; // c1t161i16
	assign leaf[233] = !f[317] && f[628] && f[545] && !f[295]; // c1t161i16
	assign leaf[234] = !f[317] && f[628] && f[545] && f[295]; // c1t161i16
	assign leaf[235] = f[317] && !f[98] && !f[99] && !f[131]; // c1t161i16
	assign leaf[236] = f[317] && !f[98] && !f[99] && f[131]; // c1t161i16
	assign leaf[237] = f[317] && !f[98] && f[99]; // c1t161i16
	assign leaf[238] = f[317] && f[98] && !f[237]; // c1t161i16
	assign leaf[239] = f[317] && f[98] && f[237]; // c1t161i16
	assign leaf[240] = !f[374] && !f[456] && !f[685] && !f[628]; // c1t171i17
	assign leaf[241] = !f[374] && !f[456] && !f[685] && f[628]; // c1t171i17
	assign leaf[242] = !f[374] && !f[456] && f[685] && !f[208]; // c1t171i17
	assign leaf[243] = !f[374] && !f[456] && f[685] && f[208]; // c1t171i17
	assign leaf[244] = !f[374] && f[456] && !f[376]; // c1t171i17
	assign leaf[245] = !f[374] && f[456] && f[376] && !f[572]; // c1t171i17
	assign leaf[246] = !f[374] && f[456] && f[376] && f[572]; // c1t171i17
	assign leaf[247] = f[374] && !f[294]; // c1t171i17
	assign leaf[248] = f[374] && f[294] && !f[126] && !f[687]; // c1t171i17
	assign leaf[249] = f[374] && f[294] && !f[126] && f[687]; // c1t171i17
	assign leaf[250] = f[374] && f[294] && f[126] && !f[491]; // c1t171i17
	assign leaf[251] = f[374] && f[294] && f[126] && f[491]; // c1t171i17
	assign leaf[252] = !f[289] && !f[351] && !f[240] && !f[184]; // c1t181i18
	assign leaf[253] = !f[289] && !f[351] && !f[240] && f[184]; // c1t181i18
	assign leaf[254] = !f[289] && !f[351] && f[240] && !f[608]; // c1t181i18
	assign leaf[255] = !f[289] && !f[351] && f[240] && f[608]; // c1t181i18
	assign leaf[256] = !f[289] && f[351] && !f[711] && !f[510]; // c1t181i18
	assign leaf[257] = !f[289] && f[351] && !f[711] && f[510]; // c1t181i18
	assign leaf[258] = !f[289] && f[351] && f[711]; // c1t181i18
	assign leaf[259] = f[289] && !f[174] && !f[98] && !f[131]; // c1t181i18
	assign leaf[260] = f[289] && !f[174] && !f[98] && f[131]; // c1t181i18
	assign leaf[261] = f[289] && !f[174] && f[98] && !f[293]; // c1t181i18
	assign leaf[262] = f[289] && !f[174] && f[98] && f[293]; // c1t181i18
	assign leaf[263] = f[289] && f[174]; // c1t181i18
	assign leaf[264] = !f[438] && !f[271] && !f[485] && !f[294]; // c1t191i19
	assign leaf[265] = !f[438] && !f[271] && !f[485] && f[294]; // c1t191i19
	assign leaf[266] = !f[438] && !f[271] && f[485] && !f[431]; // c1t191i19
	assign leaf[267] = !f[438] && !f[271] && f[485] && f[431]; // c1t191i19
	assign leaf[268] = !f[438] && f[271] && !f[183] && !f[188]; // c1t191i19
	assign leaf[269] = !f[438] && f[271] && !f[183] && f[188]; // c1t191i19
	assign leaf[270] = !f[438] && f[271] && f[183] && !f[409]; // c1t191i19
	assign leaf[271] = !f[438] && f[271] && f[183] && f[409]; // c1t191i19
	assign leaf[272] = f[438] && !f[265]; // c1t191i19
	assign leaf[273] = f[438] && f[265] && !f[152] && !f[654]; // c1t191i19
	assign leaf[274] = f[438] && f[265] && !f[152] && f[654]; // c1t191i19
	assign leaf[275] = f[438] && f[265] && f[152] && !f[491]; // c1t191i19
	assign leaf[276] = f[438] && f[265] && f[152] && f[491]; // c1t191i19
	assign leaf[277] = !f[439] && !f[683] && !f[204] && !f[537]; // c1t201i20
	assign leaf[278] = !f[439] && !f[683] && !f[204] && f[537]; // c1t201i20
	assign leaf[279] = !f[439] && !f[683] && f[204] && !f[625]; // c1t201i20
	assign leaf[280] = !f[439] && !f[683] && f[204] && f[625]; // c1t201i20
	assign leaf[281] = !f[439] && f[683] && !f[544] && !f[405]; // c1t201i20
	assign leaf[282] = !f[439] && f[683] && !f[544] && f[405]; // c1t201i20
	assign leaf[283] = !f[439] && f[683] && f[544] && !f[264]; // c1t201i20
	assign leaf[284] = !f[439] && f[683] && f[544] && f[264]; // c1t201i20
	assign leaf[285] = f[439]; // c1t201i20
	assign leaf[286] = !f[494] && !f[344] && !f[713] && !f[683]; // c1t211i21
	assign leaf[287] = !f[494] && !f[344] && !f[713] && f[683]; // c1t211i21
	assign leaf[288] = !f[494] && !f[344] && f[713] && !f[345]; // c1t211i21
	assign leaf[289] = !f[494] && !f[344] && f[713] && f[345]; // c1t211i21
	assign leaf[290] = !f[494] && f[344] && !f[128]; // c1t211i21
	assign leaf[291] = !f[494] && f[344] && f[128] && !f[153]; // c1t211i21
	assign leaf[292] = !f[494] && f[344] && f[128] && f[153]; // c1t211i21
	assign leaf[293] = f[494] && !f[125] && !f[665] && !f[72]; // c1t211i21
	assign leaf[294] = f[494] && !f[125] && !f[665] && f[72]; // c1t211i21
	assign leaf[295] = f[494] && !f[125] && f[665]; // c1t211i21
	assign leaf[296] = f[494] && f[125] && !f[237]; // c1t211i21
	assign leaf[297] = f[494] && f[125] && f[237] && !f[459]; // c1t211i21
	assign leaf[298] = f[494] && f[125] && f[237] && f[459]; // c1t211i21
	assign leaf[299] = !f[289] && !f[629] && !f[211] && !f[155]; // c1t221i22
	assign leaf[300] = !f[289] && !f[629] && !f[211] && f[155]; // c1t221i22
	assign leaf[301] = !f[289] && !f[629] && f[211] && !f[326]; // c1t221i22
	assign leaf[302] = !f[289] && !f[629] && f[211] && f[326]; // c1t221i22
	assign leaf[303] = !f[289] && f[629] && !f[545] && !f[433]; // c1t221i22
	assign leaf[304] = !f[289] && f[629] && !f[545] && f[433]; // c1t221i22
	assign leaf[305] = !f[289] && f[629] && f[545] && !f[294]; // c1t221i22
	assign leaf[306] = !f[289] && f[629] && f[545] && f[294]; // c1t221i22
	assign leaf[307] = f[289] && !f[578] && !f[606]; // c1t221i22
	assign leaf[308] = f[289] && !f[578] && f[606]; // c1t221i22
	assign leaf[309] = f[289] && f[578] && !f[491]; // c1t221i22
	assign leaf[310] = f[289] && f[578] && f[491] && !f[206]; // c1t221i22
	assign leaf[311] = f[289] && f[578] && f[491] && f[206]; // c1t221i22
	assign leaf[312] = !f[300] && !f[440] && !f[715] && !f[242]; // c1t231i23
	assign leaf[313] = !f[300] && !f[440] && !f[715] && f[242]; // c1t231i23
	assign leaf[314] = !f[300] && !f[440] && f[715] && !f[429]; // c1t231i23
	assign leaf[315] = !f[300] && !f[440] && f[715] && f[429]; // c1t231i23
	assign leaf[316] = !f[300] && f[440]; // c1t231i23
	assign leaf[317] = f[300] && !f[162] && !f[515]; // c1t231i23
	assign leaf[318] = f[300] && !f[162] && f[515] && !f[266]; // c1t231i23
	assign leaf[319] = f[300] && !f[162] && f[515] && f[266]; // c1t231i23
	assign leaf[320] = f[300] && f[162] && !f[265] && !f[573]; // c1t231i23
	assign leaf[321] = f[300] && f[162] && !f[265] && f[573]; // c1t231i23
	assign leaf[322] = f[300] && f[162] && f[265]; // c1t231i23
	assign leaf[323] = !f[711] && !f[510] && !f[344] && !f[629]; // c1t241i24
	assign leaf[324] = !f[711] && !f[510] && !f[344] && f[629]; // c1t241i24
	assign leaf[325] = !f[711] && !f[510] && f[344] && !f[597]; // c1t241i24
	assign leaf[326] = !f[711] && !f[510] && f[344] && f[597]; // c1t241i24
	assign leaf[327] = !f[711] && f[510] && !f[484]; // c1t241i24
	assign leaf[328] = !f[711] && f[510] && f[484] && !f[186]; // c1t241i24
	assign leaf[329] = !f[711] && f[510] && f[484] && f[186]; // c1t241i24
	assign leaf[330] = f[711] && !f[656]; // c1t241i24
	assign leaf[331] = f[711] && f[656] && !f[710] && !f[294]; // c1t241i24
	assign leaf[332] = f[711] && f[656] && !f[710] && f[294]; // c1t241i24
	assign leaf[333] = f[711] && f[656] && f[710] && !f[354]; // c1t241i24
	assign leaf[334] = f[711] && f[656] && f[710] && f[354]; // c1t241i24
	assign leaf[335] = !f[483] && !f[711] && !f[715] && !f[185]; // c1t251i25
	assign leaf[336] = !f[483] && !f[711] && !f[715] && f[185]; // c1t251i25
	assign leaf[337] = !f[483] && !f[711] && f[715] && !f[428]; // c1t251i25
	assign leaf[338] = !f[483] && !f[711] && f[715] && f[428]; // c1t251i25
	assign leaf[339] = !f[483] && f[711] && !f[265] && !f[460]; // c1t251i25
	assign leaf[340] = !f[483] && f[711] && !f[265] && f[460]; // c1t251i25
	assign leaf[341] = !f[483] && f[711] && f[265]; // c1t251i25
	assign leaf[342] = f[483] && !f[651] && !f[656]; // c1t251i25
	assign leaf[343] = f[483] && !f[651] && f[656] && !f[239]; // c1t251i25
	assign leaf[344] = f[483] && !f[651] && f[656] && f[239]; // c1t251i25
	assign leaf[345] = f[483] && f[651]; // c1t251i25
	assign leaf[346] = !f[209] && !f[153] && !f[265] && !f[520]; // c1t261i26
	assign leaf[347] = !f[209] && !f[153] && !f[265] && f[520]; // c1t261i26
	assign leaf[348] = !f[209] && !f[153] && f[265] && !f[155]; // c1t261i26
	assign leaf[349] = !f[209] && !f[153] && f[265] && f[155]; // c1t261i26
	assign leaf[350] = !f[209] && f[153] && !f[488] && !f[99]; // c1t261i26
	assign leaf[351] = !f[209] && f[153] && !f[488] && f[99]; // c1t261i26
	assign leaf[352] = !f[209] && f[153] && f[488] && !f[539]; // c1t261i26
	assign leaf[353] = !f[209] && f[153] && f[488] && f[539]; // c1t261i26
	assign leaf[354] = f[209] && !f[266] && !f[378] && !f[128]; // c1t261i26
	assign leaf[355] = f[209] && !f[266] && !f[378] && f[128]; // c1t261i26
	assign leaf[356] = f[209] && !f[266] && f[378] && !f[268]; // c1t261i26
	assign leaf[357] = f[209] && !f[266] && f[378] && f[268]; // c1t261i26
	assign leaf[358] = f[209] && f[266] && !f[242] && !f[177]; // c1t261i26
	assign leaf[359] = f[209] && f[266] && !f[242] && f[177]; // c1t261i26
	assign leaf[360] = f[209] && f[266] && f[242] && !f[431]; // c1t261i26
	assign leaf[361] = f[209] && f[266] && f[242] && f[431]; // c1t261i26
	assign leaf[362] = !f[383] && !f[710] && !f[492] && !f[235]; // c1t271i27
	assign leaf[363] = !f[383] && !f[710] && !f[492] && f[235]; // c1t271i27
	assign leaf[364] = !f[383] && !f[710] && f[492] && !f[606]; // c1t271i27
	assign leaf[365] = !f[383] && !f[710] && f[492] && f[606]; // c1t271i27
	assign leaf[366] = !f[383] && f[710] && !f[238] && !f[601]; // c1t271i27
	assign leaf[367] = !f[383] && f[710] && !f[238] && f[601]; // c1t271i27
	assign leaf[368] = !f[383] && f[710] && f[238]; // c1t271i27
	assign leaf[369] = f[383] && !f[218] && !f[681]; // c1t271i27
	assign leaf[370] = f[383] && !f[218] && f[681]; // c1t271i27
	assign leaf[371] = f[383] && f[218] && !f[325]; // c1t271i27
	assign leaf[372] = f[383] && f[218] && f[325]; // c1t271i27
	assign leaf[373] = !f[485] && !f[274] && !f[710] && !f[686]; // c1t281i28
	assign leaf[374] = !f[485] && !f[274] && !f[710] && f[686]; // c1t281i28
	assign leaf[375] = !f[485] && !f[274] && f[710] && !f[210]; // c1t281i28
	assign leaf[376] = !f[485] && !f[274] && f[710] && f[210]; // c1t281i28
	assign leaf[377] = !f[485] && f[274]; // c1t281i28
	assign leaf[378] = f[485] && !f[237] && !f[596] && !f[131]; // c1t281i28
	assign leaf[379] = f[485] && !f[237] && !f[596] && f[131]; // c1t281i28
	assign leaf[380] = f[485] && !f[237] && f[596] && !f[573]; // c1t281i28
	assign leaf[381] = f[485] && !f[237] && f[596] && f[573]; // c1t281i28
	assign leaf[382] = f[485] && f[237] && !f[347]; // c1t281i28
	assign leaf[383] = f[485] && f[237] && f[347] && !f[607]; // c1t281i28
	assign leaf[384] = f[485] && f[237] && f[347] && f[607]; // c1t281i28
	assign leaf[385] = !f[440] && !f[301] && !f[520] && !f[207]; // c1t291i29
	assign leaf[386] = !f[440] && !f[301] && !f[520] && f[207]; // c1t291i29
	assign leaf[387] = !f[440] && !f[301] && f[520] && !f[606]; // c1t291i29
	assign leaf[388] = !f[440] && !f[301] && f[520] && f[606]; // c1t291i29
	assign leaf[389] = !f[440] && f[301] && !f[218]; // c1t291i29
	assign leaf[390] = !f[440] && f[301] && f[218] && !f[239]; // c1t291i29
	assign leaf[391] = !f[440] && f[301] && f[218] && f[239]; // c1t291i29
	assign leaf[392] = f[440] && !f[300]; // c1t291i29
	assign leaf[393] = f[440] && f[300]; // c1t291i29
	assign leaf[394] = !f[439] && !f[272] && !f[294] && !f[182]; // c1t301i30
	assign leaf[395] = !f[439] && !f[272] && !f[294] && f[182]; // c1t301i30
	assign leaf[396] = !f[439] && !f[272] && f[294] && !f[189]; // c1t301i30
	assign leaf[397] = !f[439] && !f[272] && f[294] && f[189]; // c1t301i30
	assign leaf[398] = !f[439] && f[272] && !f[210] && !f[353]; // c1t301i30
	assign leaf[399] = !f[439] && f[272] && !f[210] && f[353]; // c1t301i30
	assign leaf[400] = !f[439] && f[272] && f[210] && !f[606]; // c1t301i30
	assign leaf[401] = !f[439] && f[272] && f[210] && f[606]; // c1t301i30
	assign leaf[402] = f[439] && !f[652]; // c1t301i30
	assign leaf[403] = f[439] && f[652]; // c1t301i30
	assign leaf[404] = !f[456] && !f[490] && !f[629] && !f[658]; // c1t311i31
	assign leaf[405] = !f[456] && !f[490] && !f[629] && f[658]; // c1t311i31
	assign leaf[406] = !f[456] && !f[490] && f[629] && !f[378]; // c1t311i31
	assign leaf[407] = !f[456] && !f[490] && f[629] && f[378]; // c1t311i31
	assign leaf[408] = !f[456] && f[490] && !f[434] && !f[580]; // c1t311i31
	assign leaf[409] = !f[456] && f[490] && !f[434] && f[580]; // c1t311i31
	assign leaf[410] = !f[456] && f[490] && f[434] && !f[244]; // c1t311i31
	assign leaf[411] = !f[456] && f[490] && f[434] && f[244]; // c1t311i31
	assign leaf[412] = f[456] && !f[658] && !f[651]; // c1t311i31
	assign leaf[413] = f[456] && !f[658] && f[651]; // c1t311i31
	assign leaf[414] = f[456] && f[658] && !f[460]; // c1t311i31
	assign leaf[415] = f[456] && f[658] && f[460]; // c1t311i31
	assign leaf[416] = !f[316] && !f[711] && !f[540] && !f[515]; // c1t321i32
	assign leaf[417] = !f[316] && !f[711] && !f[540] && f[515]; // c1t321i32
	assign leaf[418] = !f[316] && !f[711] && f[540] && !f[542]; // c1t321i32
	assign leaf[419] = !f[316] && !f[711] && f[540] && f[542]; // c1t321i32
	assign leaf[420] = !f[316] && f[711]; // c1t321i32
	assign leaf[421] = f[316] && !f[127] && !f[159] && !f[151]; // c1t321i32
	assign leaf[422] = f[316] && !f[127] && !f[159] && f[151]; // c1t321i32
	assign leaf[423] = f[316] && !f[127] && f[159]; // c1t321i32
	assign leaf[424] = f[316] && f[127] && !f[265]; // c1t321i32
	assign leaf[425] = f[316] && f[127] && f[265]; // c1t321i32
	assign leaf[426] = !f[716] && !f[713] && !f[496] && !f[185]; // c1t331i33
	assign leaf[427] = !f[716] && !f[713] && !f[496] && f[185]; // c1t331i33
	assign leaf[428] = !f[716] && !f[713] && f[496] && !f[566]; // c1t331i33
	assign leaf[429] = !f[716] && !f[713] && f[496] && f[566]; // c1t331i33
	assign leaf[430] = !f[716] && f[713] && !f[345] && !f[407]; // c1t331i33
	assign leaf[431] = !f[716] && f[713] && !f[345] && f[407]; // c1t331i33
	assign leaf[432] = !f[716] && f[713] && f[345]; // c1t331i33
	assign leaf[433] = f[716]; // c1t331i33
	assign leaf[434] = !f[537] && !f[407] && !f[463] && !f[548]; // c1t341i34
	assign leaf[435] = !f[537] && !f[407] && !f[463] && f[548]; // c1t341i34
	assign leaf[436] = !f[537] && !f[407] && f[463] && !f[460]; // c1t341i34
	assign leaf[437] = !f[537] && !f[407] && f[463] && f[460]; // c1t341i34
	assign leaf[438] = !f[537] && f[407] && !f[322] && !f[209]; // c1t341i34
	assign leaf[439] = !f[537] && f[407] && !f[322] && f[209]; // c1t341i34
	assign leaf[440] = !f[537] && f[407] && f[322] && !f[462]; // c1t341i34
	assign leaf[441] = !f[537] && f[407] && f[322] && f[462]; // c1t341i34
	assign leaf[442] = f[537] && !f[487]; // c1t341i34
	assign leaf[443] = f[537] && f[487]; // c1t341i34
	assign leaf[444] = !f[344] && !f[711] && !f[679] && !f[294]; // c1t351i35
	assign leaf[445] = !f[344] && !f[711] && !f[679] && f[294]; // c1t351i35
	assign leaf[446] = !f[344] && !f[711] && f[679] && !f[185]; // c1t351i35
	assign leaf[447] = !f[344] && !f[711] && f[679] && f[185]; // c1t351i35
	assign leaf[448] = !f[344] && f[711] && !f[710]; // c1t351i35
	assign leaf[449] = !f[344] && f[711] && f[710]; // c1t351i35
	assign leaf[450] = f[344] && !f[125] && !f[156]; // c1t351i35
	assign leaf[451] = f[344] && !f[125] && f[156] && !f[293]; // c1t351i35
	assign leaf[452] = f[344] && !f[125] && f[156] && f[293]; // c1t351i35
	assign leaf[453] = f[344] && f[125]; // c1t351i35
	assign leaf[454] = !f[440] && !f[710] && !f[407] && !f[463]; // c1t361i36
	assign leaf[455] = !f[440] && !f[710] && !f[407] && f[463]; // c1t361i36
	assign leaf[456] = !f[440] && !f[710] && f[407] && !f[578]; // c1t361i36
	assign leaf[457] = !f[440] && !f[710] && f[407] && f[578]; // c1t361i36
	assign leaf[458] = !f[440] && f[710] && !f[238]; // c1t361i36
	assign leaf[459] = !f[440] && f[710] && f[238]; // c1t361i36
	assign leaf[460] = f[440]; // c1t361i36
	assign leaf[461] = !f[511] && !f[713] && !f[537] && !f[316]; // c1t371i37
	assign leaf[462] = !f[511] && !f[713] && !f[537] && f[316]; // c1t371i37
	assign leaf[463] = !f[511] && !f[713] && f[537]; // c1t371i37
	assign leaf[464] = !f[511] && f[713] && !f[659] && !f[186]; // c1t371i37
	assign leaf[465] = !f[511] && f[713] && !f[659] && f[186]; // c1t371i37
	assign leaf[466] = !f[511] && f[713] && f[659] && !f[404]; // c1t371i37
	assign leaf[467] = !f[511] && f[713] && f[659] && f[404]; // c1t371i37
	assign leaf[468] = f[511] && !f[430] && !f[549] && !f[408]; // c1t371i37
	assign leaf[469] = f[511] && !f[430] && !f[549] && f[408]; // c1t371i37
	assign leaf[470] = f[511] && !f[430] && f[549]; // c1t371i37
	assign leaf[471] = f[511] && f[430] && !f[242]; // c1t371i37
	assign leaf[472] = f[511] && f[430] && f[242] && !f[600]; // c1t371i37
	assign leaf[473] = f[511] && f[430] && f[242] && f[600]; // c1t371i37
	assign leaf[474] = !f[621] && !f[204] && !f[565] && !f[628]; // c1t381i38
	assign leaf[475] = !f[621] && !f[204] && !f[565] && f[628]; // c1t381i38
	assign leaf[476] = !f[621] && !f[204] && f[565] && !f[488]; // c1t381i38
	assign leaf[477] = !f[621] && !f[204] && f[565] && f[488]; // c1t381i38
	assign leaf[478] = !f[621] && f[204] && !f[625] && !f[291]; // c1t381i38
	assign leaf[479] = !f[621] && f[204] && !f[625] && f[291]; // c1t381i38
	assign leaf[480] = !f[621] && f[204] && f[625] && !f[150]; // c1t381i38
	assign leaf[481] = !f[621] && f[204] && f[625] && f[150]; // c1t381i38
	assign leaf[482] = f[621] && !f[605] && !f[600] && !f[219]; // c1t381i38
	assign leaf[483] = f[621] && !f[605] && !f[600] && f[219]; // c1t381i38
	assign leaf[484] = f[621] && !f[605] && f[600]; // c1t381i38
	assign leaf[485] = f[621] && f[605]; // c1t381i38
	assign leaf[486] = !f[683] && !f[95] && !f[314] && !f[609]; // c1t391i39
	assign leaf[487] = !f[683] && !f[95] && !f[314] && f[609]; // c1t391i39
	assign leaf[488] = !f[683] && !f[95] && f[314] && !f[184]; // c1t391i39
	assign leaf[489] = !f[683] && !f[95] && f[314] && f[184]; // c1t391i39
	assign leaf[490] = !f[683] && f[95] && !f[517]; // c1t391i39
	assign leaf[491] = !f[683] && f[95] && f[517]; // c1t391i39
	assign leaf[492] = f[683] && !f[268] && !f[185]; // c1t391i39
	assign leaf[493] = f[683] && !f[268] && f[185]; // c1t391i39
	assign leaf[494] = f[683] && f[268] && !f[208] && !f[347]; // c1t391i39
	assign leaf[495] = f[683] && f[268] && !f[208] && f[347]; // c1t391i39
	assign leaf[496] = f[683] && f[268] && f[208] && !f[319]; // c1t391i39
	assign leaf[497] = f[683] && f[268] && f[208] && f[319]; // c1t391i39
	assign leaf[498] = !f[468] && !f[716] && !f[680] && !f[685]; // c1t401i40
	assign leaf[499] = !f[468] && !f[716] && !f[680] && f[685]; // c1t401i40
	assign leaf[500] = !f[468] && !f[716] && f[680] && !f[211]; // c1t401i40
	assign leaf[501] = !f[468] && !f[716] && f[680] && f[211]; // c1t401i40
	assign leaf[502] = !f[468] && f[716]; // c1t401i40
	assign leaf[503] = f[468]; // c1t401i40
	assign leaf[504] = !f[383] && !f[518] && !f[631] && !f[210]; // c1t411i41
	assign leaf[505] = !f[383] && !f[518] && !f[631] && f[210]; // c1t411i41
	assign leaf[506] = !f[383] && !f[518] && f[631] && !f[405]; // c1t411i41
	assign leaf[507] = !f[383] && !f[518] && f[631] && f[405]; // c1t411i41
	assign leaf[508] = !f[383] && f[518] && !f[603] && !f[181]; // c1t411i41
	assign leaf[509] = !f[383] && f[518] && !f[603] && f[181]; // c1t411i41
	assign leaf[510] = !f[383] && f[518] && f[603] && !f[573]; // c1t411i41
	assign leaf[511] = !f[383] && f[518] && f[603] && f[573]; // c1t411i41
	assign leaf[512] = f[383] && !f[300] && !f[380]; // c1t411i41
	assign leaf[513] = f[383] && !f[300] && f[380]; // c1t411i41
	assign leaf[514] = f[383] && f[300] && !f[213]; // c1t411i41
	assign leaf[515] = f[383] && f[300] && f[213]; // c1t411i41
	assign leaf[516] = !f[244] && !f[293] && !f[181] && !f[604]; // c1t421i42
	assign leaf[517] = !f[244] && !f[293] && !f[181] && f[604]; // c1t421i42
	assign leaf[518] = !f[244] && !f[293] && f[181] && !f[405]; // c1t421i42
	assign leaf[519] = !f[244] && !f[293] && f[181] && f[405]; // c1t421i42
	assign leaf[520] = !f[244] && f[293] && !f[160] && !f[321]; // c1t421i42
	assign leaf[521] = !f[244] && f[293] && !f[160] && f[321]; // c1t421i42
	assign leaf[522] = !f[244] && f[293] && f[160] && !f[238]; // c1t421i42
	assign leaf[523] = !f[244] && f[293] && f[160] && f[238]; // c1t421i42
	assign leaf[524] = f[244] && !f[265] && !f[156] && !f[325]; // c1t421i42
	assign leaf[525] = f[244] && !f[265] && !f[156] && f[325]; // c1t421i42
	assign leaf[526] = f[244] && !f[265] && f[156] && !f[404]; // c1t421i42
	assign leaf[527] = f[244] && !f[265] && f[156] && f[404]; // c1t421i42
	assign leaf[528] = f[244] && f[265] && !f[577] && !f[291]; // c1t421i42
	assign leaf[529] = f[244] && f[265] && !f[577] && f[291]; // c1t421i42
	assign leaf[530] = f[244] && f[265] && f[577]; // c1t421i42
	assign leaf[531] = !f[176] && !f[271] && !f[189] && !f[266]; // c1t431i43
	assign leaf[532] = !f[176] && !f[271] && !f[189] && f[266]; // c1t431i43
	assign leaf[533] = !f[176] && !f[271] && f[189] && !f[491]; // c1t431i43
	assign leaf[534] = !f[176] && !f[271] && f[189] && f[491]; // c1t431i43
	assign leaf[535] = !f[176] && f[271] && !f[381] && !f[573]; // c1t431i43
	assign leaf[536] = !f[176] && f[271] && !f[381] && f[573]; // c1t431i43
	assign leaf[537] = !f[176] && f[271] && f[381] && !f[296]; // c1t431i43
	assign leaf[538] = !f[176] && f[271] && f[381] && f[296]; // c1t431i43
	assign leaf[539] = f[176] && !f[290] && !f[127]; // c1t431i43
	assign leaf[540] = f[176] && !f[290] && f[127]; // c1t431i43
	assign leaf[541] = f[176] && f[290]; // c1t431i43
	assign leaf[542] = !f[608] && !f[260] && !f[661] && !f[292]; // c1t441i44
	assign leaf[543] = !f[608] && !f[260] && !f[661] && f[292]; // c1t441i44
	assign leaf[544] = !f[608] && !f[260] && f[661] && !f[547]; // c1t441i44
	assign leaf[545] = !f[608] && !f[260] && f[661] && f[547]; // c1t441i44
	assign leaf[546] = !f[608] && f[260] && !f[154]; // c1t441i44
	assign leaf[547] = !f[608] && f[260] && f[154]; // c1t441i44
	assign leaf[548] = f[608] && !f[488] && !f[548] && !f[625]; // c1t441i44
	assign leaf[549] = f[608] && !f[488] && !f[548] && f[625]; // c1t441i44
	assign leaf[550] = f[608] && !f[488] && f[548] && !f[267]; // c1t441i44
	assign leaf[551] = f[608] && !f[488] && f[548] && f[267]; // c1t441i44
	assign leaf[552] = f[608] && f[488] && !f[318] && !f[379]; // c1t441i44
	assign leaf[553] = f[608] && f[488] && !f[318] && f[379]; // c1t441i44
	assign leaf[554] = f[608] && f[488] && f[318]; // c1t441i44
	assign leaf[555] = !f[578] && !f[148] && !f[289] && !f[99]; // c1t451i45
	assign leaf[556] = !f[578] && !f[148] && !f[289] && f[99]; // c1t451i45
	assign leaf[557] = !f[578] && !f[148] && f[289] && !f[627]; // c1t451i45
	assign leaf[558] = !f[578] && !f[148] && f[289] && f[627]; // c1t451i45
	assign leaf[559] = !f[578] && f[148]; // c1t451i45
	assign leaf[560] = f[578] && !f[519] && !f[608] && !f[262]; // c1t451i45
	assign leaf[561] = f[578] && !f[519] && !f[608] && f[262]; // c1t451i45
	assign leaf[562] = f[578] && !f[519] && f[608] && !f[405]; // c1t451i45
	assign leaf[563] = f[578] && !f[519] && f[608] && f[405]; // c1t451i45
	assign leaf[564] = f[578] && f[519] && !f[461] && !f[350]; // c1t451i45
	assign leaf[565] = f[578] && f[519] && !f[461] && f[350]; // c1t451i45
	assign leaf[566] = f[578] && f[519] && f[461] && !f[263]; // c1t451i45
	assign leaf[567] = f[578] && f[519] && f[461] && f[263]; // c1t451i45
	assign leaf[568] = !f[578] && !f[148] && !f[493] && !f[320]; // c1t461i46
	assign leaf[569] = !f[578] && !f[148] && !f[493] && f[320]; // c1t461i46
	assign leaf[570] = !f[578] && !f[148] && f[493] && !f[237]; // c1t461i46
	assign leaf[571] = !f[578] && !f[148] && f[493] && f[237]; // c1t461i46
	assign leaf[572] = !f[578] && f[148]; // c1t461i46
	assign leaf[573] = f[578] && !f[460] && !f[491] && !f[570]; // c1t461i46
	assign leaf[574] = f[578] && !f[460] && !f[491] && f[570]; // c1t461i46
	assign leaf[575] = f[578] && !f[460] && f[491] && !f[595]; // c1t461i46
	assign leaf[576] = f[578] && !f[460] && f[491] && f[595]; // c1t461i46
	assign leaf[577] = f[578] && f[460] && !f[319] && !f[487]; // c1t461i46
	assign leaf[578] = f[578] && f[460] && !f[319] && f[487]; // c1t461i46
	assign leaf[579] = f[578] && f[460] && f[319] && !f[213]; // c1t461i46
	assign leaf[580] = f[578] && f[460] && f[319] && f[213]; // c1t461i46
	assign leaf[581] = !f[606] && !f[204] && !f[555] && !f[544]; // c1t471i47
	assign leaf[582] = !f[606] && !f[204] && !f[555] && f[544]; // c1t471i47
	assign leaf[583] = !f[606] && !f[204] && f[555]; // c1t471i47
	assign leaf[584] = !f[606] && f[204] && !f[570]; // c1t471i47
	assign leaf[585] = !f[606] && f[204] && f[570]; // c1t471i47
	assign leaf[586] = f[606] && !f[515] && !f[547] && !f[153]; // c1t471i47
	assign leaf[587] = f[606] && !f[515] && !f[547] && f[153]; // c1t471i47
	assign leaf[588] = f[606] && !f[515] && f[547] && !f[688]; // c1t471i47
	assign leaf[589] = f[606] && !f[515] && f[547] && f[688]; // c1t471i47
	assign leaf[590] = f[606] && f[515] && !f[494] && !f[431]; // c1t471i47
	assign leaf[591] = f[606] && f[515] && !f[494] && f[431]; // c1t471i47
	assign leaf[592] = f[606] && f[515] && f[494] && !f[241]; // c1t471i47
	assign leaf[593] = f[606] && f[515] && f[494] && f[241]; // c1t471i47
	assign leaf[594] = !f[271] && !f[382] && !f[459] && !f[577]; // c1t481i48
	assign leaf[595] = !f[271] && !f[382] && !f[459] && f[577]; // c1t481i48
	assign leaf[596] = !f[271] && !f[382] && f[459] && !f[377]; // c1t481i48
	assign leaf[597] = !f[271] && !f[382] && f[459] && f[377]; // c1t481i48
	assign leaf[598] = !f[271] && f[382] && !f[606] && !f[323]; // c1t481i48
	assign leaf[599] = !f[271] && f[382] && !f[606] && f[323]; // c1t481i48
	assign leaf[600] = !f[271] && f[382] && f[606]; // c1t481i48
	assign leaf[601] = f[271] && !f[408] && !f[518] && !f[157]; // c1t481i48
	assign leaf[602] = f[271] && !f[408] && !f[518] && f[157]; // c1t481i48
	assign leaf[603] = f[271] && !f[408] && f[518]; // c1t481i48
	assign leaf[604] = f[271] && f[408] && !f[132] && !f[487]; // c1t481i48
	assign leaf[605] = f[271] && f[408] && !f[132] && f[487]; // c1t481i48
	assign leaf[606] = f[271] && f[408] && f[132] && !f[156]; // c1t481i48
	assign leaf[607] = f[271] && f[408] && f[132] && f[156]; // c1t481i48
	assign leaf[608] = !f[556] && !f[260] && !f[552] && !f[99]; // c1t491i49
	assign leaf[609] = !f[556] && !f[260] && !f[552] && f[99]; // c1t491i49
	assign leaf[610] = !f[556] && !f[260] && f[552] && !f[433]; // c1t491i49
	assign leaf[611] = !f[556] && !f[260] && f[552] && f[433]; // c1t491i49
	assign leaf[612] = !f[556] && f[260] && !f[625] && !f[543]; // c1t491i49
	assign leaf[613] = !f[556] && f[260] && !f[625] && f[543]; // c1t491i49
	assign leaf[614] = !f[556] && f[260] && f[625]; // c1t491i49
	assign leaf[615] = f[556]; // c1t491i49
	assign leaf[616] = !f[96] && !f[608] && !f[510] && !f[289]; // c1t501i50
	assign leaf[617] = !f[96] && !f[608] && !f[510] && f[289]; // c1t501i50
	assign leaf[618] = !f[96] && !f[608] && f[510]; // c1t501i50
	assign leaf[619] = !f[96] && f[608] && !f[488] && !f[295]; // c1t501i50
	assign leaf[620] = !f[96] && f[608] && !f[488] && f[295]; // c1t501i50
	assign leaf[621] = !f[96] && f[608] && f[488] && !f[238]; // c1t501i50
	assign leaf[622] = !f[96] && f[608] && f[488] && f[238]; // c1t501i50
	assign leaf[623] = f[96] && !f[182]; // c1t501i50
	assign leaf[624] = f[96] && f[182]; // c1t501i50
	assign leaf[625] = !f[604] && !f[180] && !f[264] && !f[296]; // c1t511i51
	assign leaf[626] = !f[604] && !f[180] && !f[264] && f[296]; // c1t511i51
	assign leaf[627] = !f[604] && !f[180] && f[264] && !f[663]; // c1t511i51
	assign leaf[628] = !f[604] && !f[180] && f[264] && f[663]; // c1t511i51
	assign leaf[629] = !f[604] && f[180] && !f[269] && !f[125]; // c1t511i51
	assign leaf[630] = !f[604] && f[180] && !f[269] && f[125]; // c1t511i51
	assign leaf[631] = !f[604] && f[180] && f[269] && !f[152]; // c1t511i51
	assign leaf[632] = !f[604] && f[180] && f[269] && f[152]; // c1t511i51
	assign leaf[633] = f[604] && !f[546] && !f[460] && !f[658]; // c1t511i51
	assign leaf[634] = f[604] && !f[546] && !f[460] && f[658]; // c1t511i51
	assign leaf[635] = f[604] && !f[546] && f[460] && !f[576]; // c1t511i51
	assign leaf[636] = f[604] && !f[546] && f[460] && f[576]; // c1t511i51
	assign leaf[637] = f[604] && f[546] && !f[514] && !f[595]; // c1t511i51
	assign leaf[638] = f[604] && f[546] && !f[514] && f[595]; // c1t511i51
	assign leaf[639] = f[604] && f[546] && f[514] && !f[291]; // c1t511i51
	assign leaf[640] = f[604] && f[546] && f[514] && f[291]; // c1t511i51
	assign leaf[641] = !f[72] && !f[493] && !f[148] && !f[244]; // c1t521i52
	assign leaf[642] = !f[72] && !f[493] && !f[148] && f[244]; // c1t521i52
	assign leaf[643] = !f[72] && !f[493] && f[148] && !f[570]; // c1t521i52
	assign leaf[644] = !f[72] && !f[493] && f[148] && f[570]; // c1t521i52
	assign leaf[645] = !f[72] && f[493] && !f[576] && !f[179]; // c1t521i52
	assign leaf[646] = !f[72] && f[493] && !f[576] && f[179]; // c1t521i52
	assign leaf[647] = !f[72] && f[493] && f[576] && !f[519]; // c1t521i52
	assign leaf[648] = !f[72] && f[493] && f[576] && f[519]; // c1t521i52
	assign leaf[649] = f[72]; // c1t521i52
	assign leaf[650] = !f[316] && !f[627] && !f[240] && !f[185]; // c1t531i53
	assign leaf[651] = !f[316] && !f[627] && !f[240] && f[185]; // c1t531i53
	assign leaf[652] = !f[316] && !f[627] && f[240] && !f[151]; // c1t531i53
	assign leaf[653] = !f[316] && !f[627] && f[240] && f[151]; // c1t531i53
	assign leaf[654] = !f[316] && f[627] && !f[296] && !f[606]; // c1t531i53
	assign leaf[655] = !f[316] && f[627] && !f[296] && f[606]; // c1t531i53
	assign leaf[656] = !f[316] && f[627] && f[296] && !f[352]; // c1t531i53
	assign leaf[657] = !f[316] && f[627] && f[296] && f[352]; // c1t531i53
	assign leaf[658] = f[316] && !f[597]; // c1t531i53
	assign leaf[659] = f[316] && f[597]; // c1t531i53
	assign leaf[660] = !f[511] && !f[72] && !f[711] && !f[678]; // c1t541i54
	assign leaf[661] = !f[511] && !f[72] && !f[711] && f[678]; // c1t541i54
	assign leaf[662] = !f[511] && !f[72] && f[711]; // c1t541i54
	assign leaf[663] = !f[511] && f[72]; // c1t541i54
	assign leaf[664] = f[511] && !f[430] && !f[349]; // c1t541i54
	assign leaf[665] = f[511] && !f[430] && f[349]; // c1t541i54
	assign leaf[666] = f[511] && f[430] && !f[186]; // c1t541i54
	assign leaf[667] = f[511] && f[430] && f[186]; // c1t541i54
	assign leaf[668] = !f[683] && !f[411] && !f[556] && !f[606]; // c1t551i55
	assign leaf[669] = !f[683] && !f[411] && !f[556] && f[606]; // c1t551i55
	assign leaf[670] = !f[683] && !f[411] && f[556]; // c1t551i55
	assign leaf[671] = !f[683] && f[411] && !f[156]; // c1t551i55
	assign leaf[672] = !f[683] && f[411] && f[156]; // c1t551i55
	assign leaf[673] = f[683] && !f[268]; // c1t551i55
	assign leaf[674] = f[683] && f[268] && !f[207] && !f[352]; // c1t551i55
	assign leaf[675] = f[683] && f[268] && !f[207] && f[352]; // c1t551i55
	assign leaf[676] = f[683] && f[268] && f[207]; // c1t551i55
	assign leaf[677] = !f[583] && !f[152] && !f[98] && !f[236]; // c1t561i56
	assign leaf[678] = !f[583] && !f[152] && !f[98] && f[236]; // c1t561i56
	assign leaf[679] = !f[583] && !f[152] && f[98] && !f[236]; // c1t561i56
	assign leaf[680] = !f[583] && !f[152] && f[98] && f[236]; // c1t561i56
	assign leaf[681] = !f[583] && f[152] && !f[269] && !f[265]; // c1t561i56
	assign leaf[682] = !f[583] && f[152] && !f[269] && f[265]; // c1t561i56
	assign leaf[683] = !f[583] && f[152] && f[269] && !f[604]; // c1t561i56
	assign leaf[684] = !f[583] && f[152] && f[269] && f[604]; // c1t561i56
	assign leaf[685] = f[583]; // c1t561i56
	assign leaf[686] = !f[604] && !f[180] && !f[320] && !f[492]; // c1t571i57
	assign leaf[687] = !f[604] && !f[180] && !f[320] && f[492]; // c1t571i57
	assign leaf[688] = !f[604] && !f[180] && f[320] && !f[631]; // c1t571i57
	assign leaf[689] = !f[604] && !f[180] && f[320] && f[631]; // c1t571i57
	assign leaf[690] = !f[604] && f[180] && !f[269] && !f[236]; // c1t571i57
	assign leaf[691] = !f[604] && f[180] && !f[269] && f[236]; // c1t571i57
	assign leaf[692] = !f[604] && f[180] && f[269] && !f[207]; // c1t571i57
	assign leaf[693] = !f[604] && f[180] && f[269] && f[207]; // c1t571i57
	assign leaf[694] = f[604] && !f[547] && !f[266] && !f[569]; // c1t571i57
	assign leaf[695] = f[604] && !f[547] && !f[266] && f[569]; // c1t571i57
	assign leaf[696] = f[604] && !f[547] && f[266] && !f[493]; // c1t571i57
	assign leaf[697] = f[604] && !f[547] && f[266] && f[493]; // c1t571i57
	assign leaf[698] = f[604] && f[547] && !f[488] && !f[350]; // c1t571i57
	assign leaf[699] = f[604] && f[547] && !f[488] && f[350]; // c1t571i57
	assign leaf[700] = f[604] && f[547] && f[488] && !f[574]; // c1t571i57
	assign leaf[701] = f[604] && f[547] && f[488] && f[574]; // c1t571i57
	assign leaf[702] = !f[716] && !f[408] && !f[464] && !f[548]; // c1t581i58
	assign leaf[703] = !f[716] && !f[408] && !f[464] && f[548]; // c1t581i58
	assign leaf[704] = !f[716] && !f[408] && f[464] && !f[268]; // c1t581i58
	assign leaf[705] = !f[716] && !f[408] && f[464] && f[268]; // c1t581i58
	assign leaf[706] = !f[716] && f[408] && !f[324] && !f[157]; // c1t581i58
	assign leaf[707] = !f[716] && f[408] && !f[324] && f[157]; // c1t581i58
	assign leaf[708] = !f[716] && f[408] && f[324] && !f[630]; // c1t581i58
	assign leaf[709] = !f[716] && f[408] && f[324] && f[630]; // c1t581i58
	assign leaf[710] = f[716]; // c1t581i58
	assign leaf[711] = !f[609] && !f[204] && !f[157] && !f[241]; // c1t591i59
	assign leaf[712] = !f[609] && !f[204] && !f[157] && f[241]; // c1t591i59
	assign leaf[713] = !f[609] && !f[204] && f[157] && !f[268]; // c1t591i59
	assign leaf[714] = !f[609] && !f[204] && f[157] && f[268]; // c1t591i59
	assign leaf[715] = !f[609] && f[204] && !f[625] && !f[266]; // c1t591i59
	assign leaf[716] = !f[609] && f[204] && !f[625] && f[266]; // c1t591i59
	assign leaf[717] = !f[609] && f[204] && f[625]; // c1t591i59
	assign leaf[718] = f[609] && !f[157] && !f[548]; // c1t591i59
	assign leaf[719] = f[609] && !f[157] && f[548] && !f[516]; // c1t591i59
	assign leaf[720] = f[609] && !f[157] && f[548] && f[516]; // c1t591i59
	assign leaf[721] = f[609] && f[157]; // c1t591i59
	assign leaf[722] = !f[710] && !f[716] && !f[181] && !f[125]; // c1t601i60
	assign leaf[723] = !f[710] && !f[716] && !f[181] && f[125]; // c1t601i60
	assign leaf[724] = !f[710] && !f[716] && f[181] && !f[266]; // c1t601i60
	assign leaf[725] = !f[710] && !f[716] && f[181] && f[266]; // c1t601i60
	assign leaf[726] = !f[710] && f[716]; // c1t601i60
	assign leaf[727] = f[710]; // c1t601i60
	assign leaf[728] = !f[204] && !f[634] && !f[493] && !f[235]; // c1t611i61
	assign leaf[729] = !f[204] && !f[634] && !f[493] && f[235]; // c1t611i61
	assign leaf[730] = !f[204] && !f[634] && f[493] && !f[547]; // c1t611i61
	assign leaf[731] = !f[204] && !f[634] && f[493] && f[547]; // c1t611i61
	assign leaf[732] = !f[204] && f[634] && !f[348] && !f[654]; // c1t611i61
	assign leaf[733] = !f[204] && f[634] && !f[348] && f[654]; // c1t611i61
	assign leaf[734] = !f[204] && f[634] && f[348] && !f[157]; // c1t611i61
	assign leaf[735] = !f[204] && f[634] && f[348] && f[157]; // c1t611i61
	assign leaf[736] = f[204] && !f[544] && !f[599] && !f[575]; // c1t611i61
	assign leaf[737] = f[204] && !f[544] && !f[599] && f[575]; // c1t611i61
	assign leaf[738] = f[204] && !f[544] && f[599]; // c1t611i61
	assign leaf[739] = f[204] && f[544] && !f[609]; // c1t611i61
	assign leaf[740] = f[204] && f[544] && f[609]; // c1t611i61
	assign leaf[741] = !f[381] && !f[242] && !f[155] && !f[295]; // c1t621i62
	assign leaf[742] = !f[381] && !f[242] && !f[155] && f[295]; // c1t621i62
	assign leaf[743] = !f[381] && !f[242] && f[155] && !f[465]; // c1t621i62
	assign leaf[744] = !f[381] && !f[242] && f[155] && f[465]; // c1t621i62
	assign leaf[745] = !f[381] && f[242] && !f[519] && !f[183]; // c1t621i62
	assign leaf[746] = !f[381] && f[242] && !f[519] && f[183]; // c1t621i62
	assign leaf[747] = !f[381] && f[242] && f[519] && !f[408]; // c1t621i62
	assign leaf[748] = !f[381] && f[242] && f[519] && f[408]; // c1t621i62
	assign leaf[749] = f[381] && !f[297] && !f[576] && !f[460]; // c1t621i62
	assign leaf[750] = f[381] && !f[297] && !f[576] && f[460]; // c1t621i62
	assign leaf[751] = f[381] && !f[297] && f[576] && !f[125]; // c1t621i62
	assign leaf[752] = f[381] && !f[297] && f[576] && f[125]; // c1t621i62
	assign leaf[753] = f[381] && f[297] && !f[463] && !f[238]; // c1t621i62
	assign leaf[754] = f[381] && f[297] && !f[463] && f[238]; // c1t621i62
	assign leaf[755] = f[381] && f[297] && f[463] && !f[207]; // c1t621i62
	assign leaf[756] = f[381] && f[297] && f[463] && f[207]; // c1t621i62
	assign leaf[757] = !f[510] && !f[538] && !f[408] && !f[520]; // c1t631i63
	assign leaf[758] = !f[510] && !f[538] && !f[408] && f[520]; // c1t631i63
	assign leaf[759] = !f[510] && !f[538] && f[408] && !f[491]; // c1t631i63
	assign leaf[760] = !f[510] && !f[538] && f[408] && f[491]; // c1t631i63
	assign leaf[761] = !f[510] && f[538] && !f[625]; // c1t631i63
	assign leaf[762] = !f[510] && f[538] && f[625]; // c1t631i63
	assign leaf[763] = f[510]; // c1t631i63
	assign leaf[764] = !f[316] && !f[604] && !f[547] && !f[347]; // c1t641i64
	assign leaf[765] = !f[316] && !f[604] && !f[547] && f[347]; // c1t641i64
	assign leaf[766] = !f[316] && !f[604] && f[547] && !f[545]; // c1t641i64
	assign leaf[767] = !f[316] && !f[604] && f[547] && f[545]; // c1t641i64
	assign leaf[768] = !f[316] && f[604] && !f[546] && !f[460]; // c1t641i64
	assign leaf[769] = !f[316] && f[604] && !f[546] && f[460]; // c1t641i64
	assign leaf[770] = !f[316] && f[604] && f[546] && !f[102]; // c1t641i64
	assign leaf[771] = !f[316] && f[604] && f[546] && f[102]; // c1t641i64
	assign leaf[772] = f[316] && !f[126]; // c1t641i64
	assign leaf[773] = f[316] && f[126]; // c1t641i64
	assign leaf[774] = !f[102] && !f[344] && !f[132] && !f[234]; // c1t651i65
	assign leaf[775] = !f[102] && !f[344] && !f[132] && f[234]; // c1t651i65
	assign leaf[776] = !f[102] && !f[344] && f[132] && !f[520]; // c1t651i65
	assign leaf[777] = !f[102] && !f[344] && f[132] && f[520]; // c1t651i65
	assign leaf[778] = !f[102] && f[344] && !f[461]; // c1t651i65
	assign leaf[779] = !f[102] && f[344] && f[461]; // c1t651i65
	assign leaf[780] = f[102] && !f[629] && !f[626]; // c1t651i65
	assign leaf[781] = f[102] && !f[629] && f[626]; // c1t651i65
	assign leaf[782] = f[102] && f[629]; // c1t651i65
	assign leaf[783] = !f[556] && !f[511] && !f[323] && !f[183]; // c1t661i66
	assign leaf[784] = !f[556] && !f[511] && !f[323] && f[183]; // c1t661i66
	assign leaf[785] = !f[556] && !f[511] && f[323] && !f[351]; // c1t661i66
	assign leaf[786] = !f[556] && !f[511] && f[323] && f[351]; // c1t661i66
	assign leaf[787] = !f[556] && f[511] && !f[622]; // c1t661i66
	assign leaf[788] = !f[556] && f[511] && f[622]; // c1t661i66
	assign leaf[789] = f[556]; // c1t661i66
	assign leaf[790] = !f[378] && !f[322] && !f[517] && !f[434]; // c1t671i67
	assign leaf[791] = !f[378] && !f[322] && !f[517] && f[434]; // c1t671i67
	assign leaf[792] = !f[378] && !f[322] && f[517] && !f[549]; // c1t671i67
	assign leaf[793] = !f[378] && !f[322] && f[517] && f[549]; // c1t671i67
	assign leaf[794] = !f[378] && f[322] && !f[434] && !f[292]; // c1t671i67
	assign leaf[795] = !f[378] && f[322] && !f[434] && f[292]; // c1t671i67
	assign leaf[796] = !f[378] && f[322] && f[434] && !f[292]; // c1t671i67
	assign leaf[797] = !f[378] && f[322] && f[434] && f[292]; // c1t671i67
	assign leaf[798] = f[378] && !f[294] && !f[182] && !f[574]; // c1t671i67
	assign leaf[799] = f[378] && !f[294] && !f[182] && f[574]; // c1t671i67
	assign leaf[800] = f[378] && !f[294] && f[182] && !f[579]; // c1t671i67
	assign leaf[801] = f[378] && !f[294] && f[182] && f[579]; // c1t671i67
	assign leaf[802] = f[378] && f[294] && !f[375] && !f[596]; // c1t671i67
	assign leaf[803] = f[378] && f[294] && !f[375] && f[596]; // c1t671i67
	assign leaf[804] = f[378] && f[294] && f[375] && !f[657]; // c1t671i67
	assign leaf[805] = f[378] && f[294] && f[375] && f[657]; // c1t671i67
	assign leaf[806] = !f[606] && !f[204] && !f[661] && !f[263]; // c1t681i68
	assign leaf[807] = !f[606] && !f[204] && !f[661] && f[263]; // c1t681i68
	assign leaf[808] = !f[606] && !f[204] && f[661] && !f[208]; // c1t681i68
	assign leaf[809] = !f[606] && !f[204] && f[661] && f[208]; // c1t681i68
	assign leaf[810] = !f[606] && f[204] && !f[321]; // c1t681i68
	assign leaf[811] = !f[606] && f[204] && f[321]; // c1t681i68
	assign leaf[812] = f[606] && !f[267] && !f[488] && !f[547]; // c1t681i68
	assign leaf[813] = f[606] && !f[267] && !f[488] && f[547]; // c1t681i68
	assign leaf[814] = f[606] && !f[267] && f[488]; // c1t681i68
	assign leaf[815] = f[606] && f[267] && !f[149] && !f[661]; // c1t681i68
	assign leaf[816] = f[606] && f[267] && !f[149] && f[661]; // c1t681i68
	assign leaf[817] = f[606] && f[267] && f[149]; // c1t681i68
	assign leaf[818] = !f[102] && !f[213] && !f[269] && !f[321]; // c1t691i69
	assign leaf[819] = !f[102] && !f[213] && !f[269] && f[321]; // c1t691i69
	assign leaf[820] = !f[102] && !f[213] && f[269] && !f[188]; // c1t691i69
	assign leaf[821] = !f[102] && !f[213] && f[269] && f[188]; // c1t691i69
	assign leaf[822] = !f[102] && f[213] && !f[296] && !f[129]; // c1t691i69
	assign leaf[823] = !f[102] && f[213] && !f[296] && f[129]; // c1t691i69
	assign leaf[824] = !f[102] && f[213] && f[296] && !f[152]; // c1t691i69
	assign leaf[825] = !f[102] && f[213] && f[296] && f[152]; // c1t691i69
	assign leaf[826] = f[102] && !f[213]; // c1t691i69
	assign leaf[827] = f[102] && f[213]; // c1t691i69
	assign leaf[828] = !f[440] && !f[609] && !f[260] && !f[600]; // c1t701i70
	assign leaf[829] = !f[440] && !f[609] && !f[260] && f[600]; // c1t701i70
	assign leaf[830] = !f[440] && !f[609] && f[260] && !f[153]; // c1t701i70
	assign leaf[831] = !f[440] && !f[609] && f[260] && f[153]; // c1t701i70
	assign leaf[832] = !f[440] && f[609] && !f[433] && !f[157]; // c1t701i70
	assign leaf[833] = !f[440] && f[609] && !f[433] && f[157]; // c1t701i70
	assign leaf[834] = !f[440] && f[609] && f[433] && !f[376]; // c1t701i70
	assign leaf[835] = !f[440] && f[609] && f[433] && f[376]; // c1t701i70
	assign leaf[836] = f[440]; // c1t701i70
	assign leaf[837] = !f[606] && !f[289] && !f[151] && !f[99]; // c1t711i71
	assign leaf[838] = !f[606] && !f[289] && !f[151] && f[99]; // c1t711i71
	assign leaf[839] = !f[606] && !f[289] && f[151] && !f[236]; // c1t711i71
	assign leaf[840] = !f[606] && !f[289] && f[151] && f[236]; // c1t711i71
	assign leaf[841] = !f[606] && f[289]; // c1t711i71
	assign leaf[842] = f[606] && !f[491] && !f[379] && !f[461]; // c1t711i71
	assign leaf[843] = f[606] && !f[491] && !f[379] && f[461]; // c1t711i71
	assign leaf[844] = f[606] && !f[491] && f[379] && !f[626]; // c1t711i71
	assign leaf[845] = f[606] && !f[491] && f[379] && f[626]; // c1t711i71
	assign leaf[846] = f[606] && f[491] && !f[373] && !f[576]; // c1t711i71
	assign leaf[847] = f[606] && f[491] && !f[373] && f[576]; // c1t711i71
	assign leaf[848] = f[606] && f[491] && f[373]; // c1t711i71
	assign leaf[849] = !f[578] && !f[177] && !f[658] && !f[601]; // c1t721i72
	assign leaf[850] = !f[578] && !f[177] && !f[658] && f[601]; // c1t721i72
	assign leaf[851] = !f[578] && !f[177] && f[658] && !f[266]; // c1t721i72
	assign leaf[852] = !f[578] && !f[177] && f[658] && f[266]; // c1t721i72
	assign leaf[853] = !f[578] && f[177] && !f[605]; // c1t721i72
	assign leaf[854] = !f[578] && f[177] && f[605]; // c1t721i72
	assign leaf[855] = f[578] && !f[515] && !f[576] && !f[182]; // c1t721i72
	assign leaf[856] = f[578] && !f[515] && !f[576] && f[182]; // c1t721i72
	assign leaf[857] = f[578] && !f[515] && f[576] && !f[317]; // c1t721i72
	assign leaf[858] = f[578] && !f[515] && f[576] && f[317]; // c1t721i72
	assign leaf[859] = f[578] && f[515] && !f[540] && !f[375]; // c1t721i72
	assign leaf[860] = f[578] && f[515] && !f[540] && f[375]; // c1t721i72
	assign leaf[861] = f[578] && f[515] && f[540]; // c1t721i72
	assign leaf[862] = !f[381] && !f[464] && !f[324] && !f[177]; // c1t731i73
	assign leaf[863] = !f[381] && !f[464] && !f[324] && f[177]; // c1t731i73
	assign leaf[864] = !f[381] && !f[464] && f[324] && !f[264]; // c1t731i73
	assign leaf[865] = !f[381] && !f[464] && f[324] && f[264]; // c1t731i73
	assign leaf[866] = !f[381] && f[464] && !f[237] && !f[232]; // c1t731i73
	assign leaf[867] = !f[381] && f[464] && !f[237] && f[232]; // c1t731i73
	assign leaf[868] = !f[381] && f[464] && f[237] && !f[208]; // c1t731i73
	assign leaf[869] = !f[381] && f[464] && f[237] && f[208]; // c1t731i73
	assign leaf[870] = f[381] && !f[297] && !f[213] && !f[436]; // c1t731i73
	assign leaf[871] = f[381] && !f[297] && !f[213] && f[436]; // c1t731i73
	assign leaf[872] = f[381] && !f[297] && f[213] && !f[327]; // c1t731i73
	assign leaf[873] = f[381] && !f[297] && f[213] && f[327]; // c1t731i73
	assign leaf[874] = f[381] && f[297] && !f[268] && !f[595]; // c1t731i73
	assign leaf[875] = f[381] && f[297] && !f[268] && f[595]; // c1t731i73
	assign leaf[876] = f[381] && f[297] && f[268] && !f[152]; // c1t731i73
	assign leaf[877] = f[381] && f[297] && f[268] && f[152]; // c1t731i73
	assign leaf[878] = !f[555] && !f[96] && !f[378] && !f[517]; // c1t741i74
	assign leaf[879] = !f[555] && !f[96] && !f[378] && f[517]; // c1t741i74
	assign leaf[880] = !f[555] && !f[96] && f[378] && !f[322]; // c1t741i74
	assign leaf[881] = !f[555] && !f[96] && f[378] && f[322]; // c1t741i74
	assign leaf[882] = !f[555] && f[96]; // c1t741i74
	assign leaf[883] = f[555] && !f[568]; // c1t741i74
	assign leaf[884] = f[555] && f[568]; // c1t741i74
	assign leaf[885] = !f[375] && !f[321] && !f[686] && !f[460]; // c1t751i75
	assign leaf[886] = !f[375] && !f[321] && !f[686] && f[460]; // c1t751i75
	assign leaf[887] = !f[375] && !f[321] && f[686] && !f[432]; // c1t751i75
	assign leaf[888] = !f[375] && !f[321] && f[686] && f[432]; // c1t751i75
	assign leaf[889] = !f[375] && f[321] && !f[213] && !f[269]; // c1t751i75
	assign leaf[890] = !f[375] && f[321] && !f[213] && f[269]; // c1t751i75
	assign leaf[891] = !f[375] && f[321] && f[213] && !f[460]; // c1t751i75
	assign leaf[892] = !f[375] && f[321] && f[213] && f[460]; // c1t751i75
	assign leaf[893] = f[375] && !f[321] && !f[403]; // c1t751i75
	assign leaf[894] = f[375] && !f[321] && f[403]; // c1t751i75
	assign leaf[895] = f[375] && f[321] && !f[687] && !f[129]; // c1t751i75
	assign leaf[896] = f[375] && f[321] && !f[687] && f[129]; // c1t751i75
	assign leaf[897] = f[375] && f[321] && f[687] && !f[377]; // c1t751i75
	assign leaf[898] = f[375] && f[321] && f[687] && f[377]; // c1t751i75
	assign leaf[899] = !f[715] && !f[401] && !f[376] && !f[153]; // c1t761i76
	assign leaf[900] = !f[715] && !f[401] && !f[376] && f[153]; // c1t761i76
	assign leaf[901] = !f[715] && !f[401] && f[376] && !f[658]; // c1t761i76
	assign leaf[902] = !f[715] && !f[401] && f[376] && f[658]; // c1t761i76
	assign leaf[903] = !f[715] && f[401] && !f[461] && !f[345]; // c1t761i76
	assign leaf[904] = !f[715] && f[401] && !f[461] && f[345]; // c1t761i76
	assign leaf[905] = !f[715] && f[401] && f[461]; // c1t761i76
	assign leaf[906] = f[715] && !f[403]; // c1t761i76
	assign leaf[907] = f[715] && f[403]; // c1t761i76
	assign leaf[908] = !f[384] && !f[131] && !f[270] && !f[187]; // c1t771i77
	assign leaf[909] = !f[384] && !f[131] && !f[270] && f[187]; // c1t771i77
	assign leaf[910] = !f[384] && !f[131] && f[270] && !f[408]; // c1t771i77
	assign leaf[911] = !f[384] && !f[131] && f[270] && f[408]; // c1t771i77
	assign leaf[912] = !f[384] && f[131] && !f[324] && !f[129]; // c1t771i77
	assign leaf[913] = !f[384] && f[131] && !f[324] && f[129]; // c1t771i77
	assign leaf[914] = !f[384] && f[131] && f[324] && !f[241]; // c1t771i77
	assign leaf[915] = !f[384] && f[131] && f[324] && f[241]; // c1t771i77
	assign leaf[916] = f[384]; // c1t771i77
	assign leaf[917] = !f[316] && !f[635] && !f[566] && !f[540]; // c1t781i78
	assign leaf[918] = !f[316] && !f[635] && !f[566] && f[540]; // c1t781i78
	assign leaf[919] = !f[316] && !f[635] && f[566] && !f[404]; // c1t781i78
	assign leaf[920] = !f[316] && !f[635] && f[566] && f[404]; // c1t781i78
	assign leaf[921] = !f[316] && f[635] && !f[516] && !f[267]; // c1t781i78
	assign leaf[922] = !f[316] && f[635] && !f[516] && f[267]; // c1t781i78
	assign leaf[923] = !f[316] && f[635] && f[516] && !f[152]; // c1t781i78
	assign leaf[924] = !f[316] && f[635] && f[516] && f[152]; // c1t781i78
	assign leaf[925] = f[316] && !f[598]; // c1t781i78
	assign leaf[926] = f[316] && f[598]; // c1t781i78
	assign leaf[927] = !f[603] && !f[209] && !f[265] && !f[346]; // c1t791i79
	assign leaf[928] = !f[603] && !f[209] && !f[265] && f[346]; // c1t791i79
	assign leaf[929] = !f[603] && !f[209] && f[265] && !f[636]; // c1t791i79
	assign leaf[930] = !f[603] && !f[209] && f[265] && f[636]; // c1t791i79
	assign leaf[931] = !f[603] && f[209] && !f[238] && !f[295]; // c1t791i79
	assign leaf[932] = !f[603] && f[209] && !f[238] && f[295]; // c1t791i79
	assign leaf[933] = !f[603] && f[209] && f[238] && !f[325]; // c1t791i79
	assign leaf[934] = !f[603] && f[209] && f[238] && f[325]; // c1t791i79
	assign leaf[935] = f[603] && !f[546] && !f[578] && !f[210]; // c1t791i79
	assign leaf[936] = f[603] && !f[546] && !f[578] && f[210]; // c1t791i79
	assign leaf[937] = f[603] && !f[546] && f[578] && !f[492]; // c1t791i79
	assign leaf[938] = f[603] && !f[546] && f[578] && f[492]; // c1t791i79
	assign leaf[939] = f[603] && f[546] && !f[241] && !f[158]; // c1t791i79
	assign leaf[940] = f[603] && f[546] && !f[241] && f[158]; // c1t791i79
	assign leaf[941] = f[603] && f[546] && f[241] && !f[129]; // c1t791i79
	assign leaf[942] = f[603] && f[546] && f[241] && f[129]; // c1t791i79
	assign leaf[943] = !f[440] && !f[204] && !f[658] && !f[517]; // c1t801i80
	assign leaf[944] = !f[440] && !f[204] && !f[658] && f[517]; // c1t801i80
	assign leaf[945] = !f[440] && !f[204] && f[658] && !f[436]; // c1t801i80
	assign leaf[946] = !f[440] && !f[204] && f[658] && f[436]; // c1t801i80
	assign leaf[947] = !f[440] && f[204] && !f[291] && !f[269]; // c1t801i80
	assign leaf[948] = !f[440] && f[204] && !f[291] && f[269]; // c1t801i80
	assign leaf[949] = !f[440] && f[204] && f[291]; // c1t801i80
	assign leaf[950] = f[440]; // c1t801i80
	assign leaf[951] = !f[456] && !f[686] && !f[578] && !f[433]; // c1t811i81
	assign leaf[952] = !f[456] && !f[686] && !f[578] && f[433]; // c1t811i81
	assign leaf[953] = !f[456] && !f[686] && f[578] && !f[491]; // c1t811i81
	assign leaf[954] = !f[456] && !f[686] && f[578] && f[491]; // c1t811i81
	assign leaf[955] = !f[456] && f[686] && !f[180] && !f[263]; // c1t811i81
	assign leaf[956] = !f[456] && f[686] && !f[180] && f[263]; // c1t811i81
	assign leaf[957] = !f[456] && f[686] && f[180] && !f[347]; // c1t811i81
	assign leaf[958] = !f[456] && f[686] && f[180] && f[347]; // c1t811i81
	assign leaf[959] = f[456] && !f[630]; // c1t811i81
	assign leaf[960] = f[456] && f[630]; // c1t811i81
	assign leaf[961] = !f[329] && !f[375] && !f[321] && !f[181]; // c1t821i82
	assign leaf[962] = !f[329] && !f[375] && !f[321] && f[181]; // c1t821i82
	assign leaf[963] = !f[329] && !f[375] && f[321] && !f[622]; // c1t821i82
	assign leaf[964] = !f[329] && !f[375] && f[321] && f[622]; // c1t821i82
	assign leaf[965] = !f[329] && f[375] && !f[321] && !f[548]; // c1t821i82
	assign leaf[966] = !f[329] && f[375] && !f[321] && f[548]; // c1t821i82
	assign leaf[967] = !f[329] && f[375] && f[321] && !f[658]; // c1t821i82
	assign leaf[968] = !f[329] && f[375] && f[321] && f[658]; // c1t821i82
	assign leaf[969] = f[329]; // c1t821i82
	assign leaf[970] = !f[709] && !f[204] && !f[245] && !f[538]; // c1t831i83
	assign leaf[971] = !f[709] && !f[204] && !f[245] && f[538]; // c1t831i83
	assign leaf[972] = !f[709] && !f[204] && f[245] && !f[162]; // c1t831i83
	assign leaf[973] = !f[709] && !f[204] && f[245] && f[162]; // c1t831i83
	assign leaf[974] = !f[709] && f[204] && !f[569] && !f[636]; // c1t831i83
	assign leaf[975] = !f[709] && f[204] && !f[569] && f[636]; // c1t831i83
	assign leaf[976] = !f[709] && f[204] && f[569]; // c1t831i83
	assign leaf[977] = f[709]; // c1t831i83
	assign leaf[978] = !f[708] && !f[244] && !f[204] && !f[266]; // c1t841i84
	assign leaf[979] = !f[708] && !f[244] && !f[204] && f[266]; // c1t841i84
	assign leaf[980] = !f[708] && !f[244] && f[204] && !f[156]; // c1t841i84
	assign leaf[981] = !f[708] && !f[244] && f[204] && f[156]; // c1t841i84
	assign leaf[982] = !f[708] && f[244] && !f[293] && !f[129]; // c1t841i84
	assign leaf[983] = !f[708] && f[244] && !f[293] && f[129]; // c1t841i84
	assign leaf[984] = !f[708] && f[244] && f[293] && !f[595]; // c1t841i84
	assign leaf[985] = !f[708] && f[244] && f[293] && f[595]; // c1t841i84
	assign leaf[986] = f[708]; // c1t841i84
	assign leaf[987] = !f[493] && !f[519] && !f[464] && !f[353]; // c1t851i85
	assign leaf[988] = !f[493] && !f[519] && !f[464] && f[353]; // c1t851i85
	assign leaf[989] = !f[493] && !f[519] && f[464] && !f[487]; // c1t851i85
	assign leaf[990] = !f[493] && !f[519] && f[464] && f[487]; // c1t851i85
	assign leaf[991] = !f[493] && f[519] && !f[546] && !f[180]; // c1t851i85
	assign leaf[992] = !f[493] && f[519] && !f[546] && f[180]; // c1t851i85
	assign leaf[993] = !f[493] && f[519] && f[546] && !f[462]; // c1t851i85
	assign leaf[994] = !f[493] && f[519] && f[546] && f[462]; // c1t851i85
	assign leaf[995] = f[493] && !f[636] && !f[547]; // c1t851i85
	assign leaf[996] = f[493] && !f[636] && f[547] && !f[265]; // c1t851i85
	assign leaf[997] = f[493] && !f[636] && f[547] && f[265]; // c1t851i85
	assign leaf[998] = f[493] && f[636]; // c1t851i85
	assign leaf[999] = !f[356] && !f[215] && !f[353] && !f[566]; // c1t861i86
	assign leaf[1000] = !f[356] && !f[215] && !f[353] && f[566]; // c1t861i86
	assign leaf[1001] = !f[356] && !f[215] && f[353] && !f[659]; // c1t861i86
	assign leaf[1002] = !f[356] && !f[215] && f[353] && f[659]; // c1t861i86
	assign leaf[1003] = !f[356] && f[215] && !f[381] && !f[519]; // c1t861i86
	assign leaf[1004] = !f[356] && f[215] && !f[381] && f[519]; // c1t861i86
	assign leaf[1005] = !f[356] && f[215] && f[381] && !f[436]; // c1t861i86
	assign leaf[1006] = !f[356] && f[215] && f[381] && f[436]; // c1t861i86
	assign leaf[1007] = f[356]; // c1t861i86
	assign leaf[1008] = !f[152] && !f[656] && !f[573] && !f[714]; // c1t871i87
	assign leaf[1009] = !f[152] && !f[656] && !f[573] && f[714]; // c1t871i87
	assign leaf[1010] = !f[152] && !f[656] && f[573] && !f[486]; // c1t871i87
	assign leaf[1011] = !f[152] && !f[656] && f[573] && f[486]; // c1t871i87
	assign leaf[1012] = !f[152] && f[656] && !f[380] && !f[270]; // c1t871i87
	assign leaf[1013] = !f[152] && f[656] && !f[380] && f[270]; // c1t871i87
	assign leaf[1014] = !f[152] && f[656] && f[380] && !f[463]; // c1t871i87
	assign leaf[1015] = !f[152] && f[656] && f[380] && f[463]; // c1t871i87
	assign leaf[1016] = f[152] && !f[269] && !f[236] && !f[206]; // c1t871i87
	assign leaf[1017] = f[152] && !f[269] && !f[236] && f[206]; // c1t871i87
	assign leaf[1018] = f[152] && !f[269] && f[236] && !f[547]; // c1t871i87
	assign leaf[1019] = f[152] && !f[269] && f[236] && f[547]; // c1t871i87
	assign leaf[1020] = f[152] && f[269] && !f[462]; // c1t871i87
	assign leaf[1021] = f[152] && f[269] && f[462] && !f[375]; // c1t871i87
	assign leaf[1022] = f[152] && f[269] && f[462] && f[375]; // c1t871i87
	assign leaf[1023] = !f[244] && !f[566] && !f[493] && !f[178]; // c1t881i88
	assign leaf[1024] = !f[244] && !f[566] && !f[493] && f[178]; // c1t881i88
	assign leaf[1025] = !f[244] && !f[566] && f[493] && !f[519]; // c1t881i88
	assign leaf[1026] = !f[244] && !f[566] && f[493] && f[519]; // c1t881i88
	assign leaf[1027] = !f[244] && f[566] && !f[349]; // c1t881i88
	assign leaf[1028] = !f[244] && f[566] && f[349]; // c1t881i88
	assign leaf[1029] = f[244] && !f[321] && !f[381]; // c1t881i88
	assign leaf[1030] = f[244] && !f[321] && f[381] && !f[296]; // c1t881i88
	assign leaf[1031] = f[244] && !f[321] && f[381] && f[296]; // c1t881i88
	assign leaf[1032] = f[244] && f[321] && !f[320] && !f[430]; // c1t881i88
	assign leaf[1033] = f[244] && f[321] && !f[320] && f[430]; // c1t881i88
	assign leaf[1034] = f[244] && f[321] && f[320]; // c1t881i88
	assign leaf[1035] = !f[713] && !f[548] && !f[151] && !f[569]; // c1t891i89
	assign leaf[1036] = !f[713] && !f[548] && !f[151] && f[569]; // c1t891i89
	assign leaf[1037] = !f[713] && !f[548] && f[151] && !f[659]; // c1t891i89
	assign leaf[1038] = !f[713] && !f[548] && f[151] && f[659]; // c1t891i89
	assign leaf[1039] = !f[713] && f[548] && !f[576] && !f[129]; // c1t891i89
	assign leaf[1040] = !f[713] && f[548] && !f[576] && f[129]; // c1t891i89
	assign leaf[1041] = !f[713] && f[548] && f[576] && !f[405]; // c1t891i89
	assign leaf[1042] = !f[713] && f[548] && f[576] && f[405]; // c1t891i89
	assign leaf[1043] = f[713] && !f[349]; // c1t891i89
	assign leaf[1044] = f[713] && f[349]; // c1t891i89
	assign leaf[1045] = !f[712] && !f[440] && !f[578] && !f[177]; // c1t901i90
	assign leaf[1046] = !f[712] && !f[440] && !f[578] && f[177]; // c1t901i90
	assign leaf[1047] = !f[712] && !f[440] && f[578] && !f[517]; // c1t901i90
	assign leaf[1048] = !f[712] && !f[440] && f[578] && f[517]; // c1t901i90
	assign leaf[1049] = !f[712] && f[440]; // c1t901i90
	assign leaf[1050] = f[712] && !f[432]; // c1t901i90
	assign leaf[1051] = f[712] && f[432]; // c1t901i90
	assign leaf[1052] = !f[215] && !f[381] && !f[241] && !f[210]; // c1t911i91
	assign leaf[1053] = !f[215] && !f[381] && !f[241] && f[210]; // c1t911i91
	assign leaf[1054] = !f[215] && !f[381] && f[241] && !f[575]; // c1t911i91
	assign leaf[1055] = !f[215] && !f[381] && f[241] && f[575]; // c1t911i91
	assign leaf[1056] = !f[215] && f[381] && !f[548] && !f[240]; // c1t911i91
	assign leaf[1057] = !f[215] && f[381] && !f[548] && f[240]; // c1t911i91
	assign leaf[1058] = !f[215] && f[381] && f[548] && !f[346]; // c1t911i91
	assign leaf[1059] = !f[215] && f[381] && f[548] && f[346]; // c1t911i91
	assign leaf[1060] = f[215] && !f[324]; // c1t911i91
	assign leaf[1061] = f[215] && f[324] && !f[381] && !f[519]; // c1t911i91
	assign leaf[1062] = f[215] && f[324] && !f[381] && f[519]; // c1t911i91
	assign leaf[1063] = f[215] && f[324] && f[381] && !f[209]; // c1t911i91
	assign leaf[1064] = f[215] && f[324] && f[381] && f[209]; // c1t911i91
	assign leaf[1065] = !f[95] && !f[609] && !f[708] && !f[204]; // c1t921i92
	assign leaf[1066] = !f[95] && !f[609] && !f[708] && f[204]; // c1t921i92
	assign leaf[1067] = !f[95] && !f[609] && f[708]; // c1t921i92
	assign leaf[1068] = !f[95] && f[609] && !f[516]; // c1t921i92
	assign leaf[1069] = !f[95] && f[609] && f[516]; // c1t921i92
	assign leaf[1070] = f[95]; // c1t921i92
	assign leaf[1071] = !f[715] && !f[712] && !f[374] && !f[244]; // c1t931i93
	assign leaf[1072] = !f[715] && !f[712] && !f[374] && f[244]; // c1t931i93
	assign leaf[1073] = !f[715] && !f[712] && f[374] && !f[323]; // c1t931i93
	assign leaf[1074] = !f[715] && !f[712] && f[374] && f[323]; // c1t931i93
	assign leaf[1075] = !f[715] && f[712] && !f[376]; // c1t931i93
	assign leaf[1076] = !f[715] && f[712] && f[376]; // c1t931i93
	assign leaf[1077] = f[715] && !f[346]; // c1t931i93
	assign leaf[1078] = f[715] && f[346]; // c1t931i93
	assign leaf[1079] = !f[490] && !f[378] && !f[322] && !f[434]; // c1t941i94
	assign leaf[1080] = !f[490] && !f[378] && !f[322] && f[434]; // c1t941i94
	assign leaf[1081] = !f[490] && !f[378] && f[322]; // c1t941i94
	assign leaf[1082] = !f[490] && f[378] && !f[630] && !f[569]; // c1t941i94
	assign leaf[1083] = !f[490] && f[378] && !f[630] && f[569]; // c1t941i94
	assign leaf[1084] = !f[490] && f[378] && f[630] && !f[407]; // c1t941i94
	assign leaf[1085] = !f[490] && f[378] && f[630] && f[407]; // c1t941i94
	assign leaf[1086] = f[490] && !f[603] && !f[516] && !f[635]; // c1t941i94
	assign leaf[1087] = f[490] && !f[603] && !f[516] && f[635]; // c1t941i94
	assign leaf[1088] = f[490] && !f[603] && f[516] && !f[236]; // c1t941i94
	assign leaf[1089] = f[490] && !f[603] && f[516] && f[236]; // c1t941i94
	assign leaf[1090] = f[490] && f[603] && !f[573] && !f[488]; // c1t941i94
	assign leaf[1091] = f[490] && f[603] && !f[573] && f[488]; // c1t941i94
	assign leaf[1092] = f[490] && f[603] && f[573] && !f[177]; // c1t941i94
	assign leaf[1093] = f[490] && f[603] && f[573] && f[177]; // c1t941i94
	assign leaf[1094] = !f[378] && !f[682] && !f[624] && !f[321]; // c1t951i95
	assign leaf[1095] = !f[378] && !f[682] && !f[624] && f[321]; // c1t951i95
	assign leaf[1096] = !f[378] && !f[682] && f[624] && !f[379]; // c1t951i95
	assign leaf[1097] = !f[378] && !f[682] && f[624] && f[379]; // c1t951i95
	assign leaf[1098] = !f[378] && f[682]; // c1t951i95
	assign leaf[1099] = f[378] && !f[294] && !f[539] && !f[403]; // c1t951i95
	assign leaf[1100] = f[378] && !f[294] && !f[539] && f[403]; // c1t951i95
	assign leaf[1101] = f[378] && !f[294] && f[539]; // c1t951i95
	assign leaf[1102] = f[378] && f[294] && !f[322]; // c1t951i95
	assign leaf[1103] = f[378] && f[294] && f[322] && !f[177]; // c1t951i95
	assign leaf[1104] = f[378] && f[294] && f[322] && f[177]; // c1t951i95
	assign leaf[1105] = !f[265] && !f[155] && !f[241] && !f[295]; // c1t961i96
	assign leaf[1106] = !f[265] && !f[155] && !f[241] && f[295]; // c1t961i96
	assign leaf[1107] = !f[265] && !f[155] && f[241] && !f[324]; // c1t961i96
	assign leaf[1108] = !f[265] && !f[155] && f[241] && f[324]; // c1t961i96
	assign leaf[1109] = !f[265] && f[155] && !f[239] && !f[406]; // c1t961i96
	assign leaf[1110] = !f[265] && f[155] && !f[239] && f[406]; // c1t961i96
	assign leaf[1111] = !f[265] && f[155] && f[239] && !f[487]; // c1t961i96
	assign leaf[1112] = !f[265] && f[155] && f[239] && f[487]; // c1t961i96
	assign leaf[1113] = f[265] && !f[159] && !f[349] && !f[157]; // c1t961i96
	assign leaf[1114] = f[265] && !f[159] && !f[349] && f[157]; // c1t961i96
	assign leaf[1115] = f[265] && !f[159] && f[349] && !f[431]; // c1t961i96
	assign leaf[1116] = f[265] && !f[159] && f[349] && f[431]; // c1t961i96
	assign leaf[1117] = f[265] && f[159] && !f[406]; // c1t961i96
	assign leaf[1118] = f[265] && f[159] && f[406] && !f[486]; // c1t961i96
	assign leaf[1119] = f[265] && f[159] && f[406] && f[486]; // c1t961i96
	assign leaf[1120] = !f[658] && !f[517] && !f[184] && !f[238]; // c1t971i97
	assign leaf[1121] = !f[658] && !f[517] && !f[184] && f[238]; // c1t971i97
	assign leaf[1122] = !f[658] && !f[517] && f[184] && !f[578]; // c1t971i97
	assign leaf[1123] = !f[658] && !f[517] && f[184] && f[578]; // c1t971i97
	assign leaf[1124] = !f[658] && f[517] && !f[241] && !f[380]; // c1t971i97
	assign leaf[1125] = !f[658] && f[517] && !f[241] && f[380]; // c1t971i97
	assign leaf[1126] = !f[658] && f[517] && f[241] && !f[349]; // c1t971i97
	assign leaf[1127] = !f[658] && f[517] && f[241] && f[349]; // c1t971i97
	assign leaf[1128] = f[658] && !f[266] && !f[181]; // c1t971i97
	assign leaf[1129] = f[658] && !f[266] && f[181] && !f[464]; // c1t971i97
	assign leaf[1130] = f[658] && !f[266] && f[181] && f[464]; // c1t971i97
	assign leaf[1131] = f[658] && f[266] && !f[517] && !f[377]; // c1t971i97
	assign leaf[1132] = f[658] && f[266] && !f[517] && f[377]; // c1t971i97
	assign leaf[1133] = f[658] && f[266] && f[517] && !f[600]; // c1t971i97
	assign leaf[1134] = f[658] && f[266] && f[517] && f[600]; // c1t971i97
	assign leaf[1135] = !f[320] && !f[687] && !f[373] && !f[657]; // c1t981i98
	assign leaf[1136] = !f[320] && !f[687] && !f[373] && f[657]; // c1t981i98
	assign leaf[1137] = !f[320] && !f[687] && f[373]; // c1t981i98
	assign leaf[1138] = !f[320] && f[687] && !f[180]; // c1t981i98
	assign leaf[1139] = !f[320] && f[687] && f[180] && !f[154]; // c1t981i98
	assign leaf[1140] = !f[320] && f[687] && f[180] && f[154]; // c1t981i98
	assign leaf[1141] = f[320] && !f[662] && !f[460] && !f[547]; // c1t981i98
	assign leaf[1142] = f[320] && !f[662] && !f[460] && f[547]; // c1t981i98
	assign leaf[1143] = f[320] && !f[662] && f[460] && !f[405]; // c1t981i98
	assign leaf[1144] = f[320] && !f[662] && f[460] && f[405]; // c1t981i98
	assign leaf[1145] = f[320] && f[662] && !f[267]; // c1t981i98
	assign leaf[1146] = f[320] && f[662] && f[267]; // c1t981i98
	assign leaf[1147] = !f[708] && !f[403] && !f[714] && !f[321]; // c1t991i99
	assign leaf[1148] = !f[708] && !f[403] && !f[714] && f[321]; // c1t991i99
	assign leaf[1149] = !f[708] && !f[403] && f[714] && !f[184]; // c1t991i99
	assign leaf[1150] = !f[708] && !f[403] && f[714] && f[184]; // c1t991i99
	assign leaf[1151] = !f[708] && f[403] && !f[349]; // c1t991i99
	assign leaf[1152] = !f[708] && f[403] && f[349] && !f[155]; // c1t991i99
	assign leaf[1153] = !f[708] && f[403] && f[349] && f[155]; // c1t991i99
	assign leaf[1154] = f[708]; // c1t991i99
endmodule

module decision_tree_leaves_2(input logic [0:783] f, output logic [0:1374] leaf);
	assign leaf[0] = !f[583] && !f[124] && !f[528] && !f[564]; // c2t2i0
	assign leaf[1] = !f[583] && !f[124] && !f[528] && f[564]; // c2t2i0
	assign leaf[2] = !f[583] && !f[124] && f[528] && !f[371]; // c2t2i0
	assign leaf[3] = !f[583] && !f[124] && f[528] && f[371]; // c2t2i0
	assign leaf[4] = !f[583] && f[124] && !f[346] && !f[349]; // c2t2i0
	assign leaf[5] = !f[583] && f[124] && !f[346] && f[349]; // c2t2i0
	assign leaf[6] = !f[583] && f[124] && f[346] && !f[93]; // c2t2i0
	assign leaf[7] = !f[583] && f[124] && f[346] && f[93]; // c2t2i0
	assign leaf[8] = f[583] && !f[343] && !f[346] && !f[369]; // c2t2i0
	assign leaf[9] = f[583] && !f[343] && !f[346] && f[369]; // c2t2i0
	assign leaf[10] = f[583] && !f[343] && f[346] && !f[520]; // c2t2i0
	assign leaf[11] = f[583] && !f[343] && f[346] && f[520]; // c2t2i0
	assign leaf[12] = f[583] && f[343] && !f[519] && !f[517]; // c2t2i0
	assign leaf[13] = f[583] && f[343] && !f[519] && f[517]; // c2t2i0
	assign leaf[14] = f[583] && f[343] && f[519] && !f[442]; // c2t2i0
	assign leaf[15] = f[583] && f[343] && f[519] && f[442]; // c2t2i0
	assign leaf[16] = !f[542] && !f[512] && !f[99] && !f[571]; // c2t12i1
	assign leaf[17] = !f[542] && !f[512] && !f[99] && f[571]; // c2t12i1
	assign leaf[18] = !f[542] && !f[512] && f[99] && !f[482]; // c2t12i1
	assign leaf[19] = !f[542] && !f[512] && f[99] && f[482]; // c2t12i1
	assign leaf[20] = !f[542] && f[512] && !f[346] && !f[658]; // c2t12i1
	assign leaf[21] = !f[542] && f[512] && !f[346] && f[658]; // c2t12i1
	assign leaf[22] = !f[542] && f[512] && f[346] && !f[97]; // c2t12i1
	assign leaf[23] = !f[542] && f[512] && f[346] && f[97]; // c2t12i1
	assign leaf[24] = f[542] && !f[347] && !f[344] && !f[350]; // c2t12i1
	assign leaf[25] = f[542] && !f[347] && !f[344] && f[350]; // c2t12i1
	assign leaf[26] = f[542] && !f[347] && f[344] && !f[372]; // c2t12i1
	assign leaf[27] = f[542] && !f[347] && f[344] && f[372]; // c2t12i1
	assign leaf[28] = f[542] && f[347] && !f[528] && !f[582]; // c2t12i1
	assign leaf[29] = f[542] && f[347] && !f[528] && f[582]; // c2t12i1
	assign leaf[30] = f[542] && f[347] && f[528] && !f[414]; // c2t12i1
	assign leaf[31] = f[542] && f[347] && f[528] && f[414]; // c2t12i1
	assign leaf[32] = !f[568] && !f[123] && !f[539] && !f[473]; // c2t22i2
	assign leaf[33] = !f[568] && !f[123] && !f[539] && f[473]; // c2t22i2
	assign leaf[34] = !f[568] && !f[123] && f[539] && !f[346]; // c2t22i2
	assign leaf[35] = !f[568] && !f[123] && f[539] && f[346]; // c2t22i2
	assign leaf[36] = !f[568] && f[123] && !f[345] && !f[348]; // c2t22i2
	assign leaf[37] = !f[568] && f[123] && !f[345] && f[348]; // c2t22i2
	assign leaf[38] = !f[568] && f[123] && f[345] && !f[664]; // c2t22i2
	assign leaf[39] = !f[568] && f[123] && f[345] && f[664]; // c2t22i2
	assign leaf[40] = f[568] && !f[517] && !f[460] && !f[98]; // c2t22i2
	assign leaf[41] = f[568] && !f[517] && !f[460] && f[98]; // c2t22i2
	assign leaf[42] = f[568] && !f[517] && f[460] && !f[348]; // c2t22i2
	assign leaf[43] = f[568] && !f[517] && f[460] && f[348]; // c2t22i2
	assign leaf[44] = f[568] && f[517] && !f[320] && !f[156]; // c2t22i2
	assign leaf[45] = f[568] && f[517] && !f[320] && f[156]; // c2t22i2
	assign leaf[46] = f[568] && f[517] && f[320] && !f[580]; // c2t22i2
	assign leaf[47] = f[568] && f[517] && f[320] && f[580]; // c2t22i2
	assign leaf[48] = !f[346] && !f[569] && !f[511] && !f[582]; // c2t32i3
	assign leaf[49] = !f[346] && !f[569] && !f[511] && f[582]; // c2t32i3
	assign leaf[50] = !f[346] && !f[569] && f[511] && !f[343]; // c2t32i3
	assign leaf[51] = !f[346] && !f[569] && f[511] && f[343]; // c2t32i3
	assign leaf[52] = !f[346] && f[569] && !f[321] && !f[371]; // c2t32i3
	assign leaf[53] = !f[346] && f[569] && !f[321] && f[371]; // c2t32i3
	assign leaf[54] = !f[346] && f[569] && f[321] && !f[554]; // c2t32i3
	assign leaf[55] = !f[346] && f[569] && f[321] && f[554]; // c2t32i3
	assign leaf[56] = f[346] && !f[528] && !f[584] && !f[637]; // c2t32i3
	assign leaf[57] = f[346] && !f[528] && !f[584] && f[637]; // c2t32i3
	assign leaf[58] = f[346] && !f[528] && f[584]; // c2t32i3
	assign leaf[59] = f[346] && f[528] && !f[413] && !f[551]; // c2t32i3
	assign leaf[60] = f[346] && f[528] && !f[413] && f[551]; // c2t32i3
	assign leaf[61] = f[346] && f[528] && f[413] && !f[493]; // c2t32i3
	assign leaf[62] = f[346] && f[528] && f[413] && f[493]; // c2t32i3
	assign leaf[63] = !f[345] && !f[348] && !f[153] && !f[538]; // c2t42i4
	assign leaf[64] = !f[345] && !f[348] && !f[153] && f[538]; // c2t42i4
	assign leaf[65] = !f[345] && !f[348] && f[153] && !f[516]; // c2t42i4
	assign leaf[66] = !f[345] && !f[348] && f[153] && f[516]; // c2t42i4
	assign leaf[67] = !f[345] && f[348] && !f[473] && !f[554]; // c2t42i4
	assign leaf[68] = !f[345] && f[348] && !f[473] && f[554]; // c2t42i4
	assign leaf[69] = !f[345] && f[348] && f[473] && !f[528]; // c2t42i4
	assign leaf[70] = !f[345] && f[348] && f[473] && f[528]; // c2t42i4
	assign leaf[71] = f[345] && !f[583] && !f[501] && !f[568]; // c2t42i4
	assign leaf[72] = f[345] && !f[583] && !f[501] && f[568]; // c2t42i4
	assign leaf[73] = f[345] && !f[583] && f[501] && !f[267]; // c2t42i4
	assign leaf[74] = f[345] && !f[583] && f[501] && f[267]; // c2t42i4
	assign leaf[75] = f[345] && f[583] && !f[518] && !f[490]; // c2t42i4
	assign leaf[76] = f[345] && f[583] && !f[518] && f[490]; // c2t42i4
	assign leaf[77] = f[345] && f[583] && f[518] && !f[430]; // c2t42i4
	assign leaf[78] = f[345] && f[583] && f[518] && f[430]; // c2t42i4
	assign leaf[79] = !f[543] && !f[512] && !f[99] && !f[514]; // c2t52i5
	assign leaf[80] = !f[543] && !f[512] && !f[99] && f[514]; // c2t52i5
	assign leaf[81] = !f[543] && !f[512] && f[99] && !f[351]; // c2t52i5
	assign leaf[82] = !f[543] && !f[512] && f[99] && f[351]; // c2t52i5
	assign leaf[83] = !f[543] && f[512] && !f[319] && !f[316]; // c2t52i5
	assign leaf[84] = !f[543] && f[512] && !f[319] && f[316]; // c2t52i5
	assign leaf[85] = !f[543] && f[512] && f[319] && !f[630]; // c2t52i5
	assign leaf[86] = !f[543] && f[512] && f[319] && f[630]; // c2t52i5
	assign leaf[87] = f[543] && !f[346] && !f[181] && !f[126]; // c2t52i5
	assign leaf[88] = f[543] && !f[346] && !f[181] && f[126]; // c2t52i5
	assign leaf[89] = f[543] && !f[346] && f[181] && !f[371]; // c2t52i5
	assign leaf[90] = f[543] && !f[346] && f[181] && f[371]; // c2t52i5
	assign leaf[91] = f[543] && f[346] && !f[318] && !f[426]; // c2t52i5
	assign leaf[92] = f[543] && f[346] && !f[318] && f[426]; // c2t52i5
	assign leaf[93] = f[543] && f[346] && f[318] && !f[374]; // c2t52i5
	assign leaf[94] = f[543] && f[346] && f[318] && f[374]; // c2t52i5
	assign leaf[95] = !f[346] && !f[543] && !f[485] && !f[514]; // c2t62i6
	assign leaf[96] = !f[346] && !f[543] && !f[485] && f[514]; // c2t62i6
	assign leaf[97] = !f[346] && !f[543] && f[485] && !f[343]; // c2t62i6
	assign leaf[98] = !f[346] && !f[543] && f[485] && f[343]; // c2t62i6
	assign leaf[99] = !f[346] && f[543] && !f[154] && !f[653]; // c2t62i6
	assign leaf[100] = !f[346] && f[543] && !f[154] && f[653]; // c2t62i6
	assign leaf[101] = !f[346] && f[543] && f[154] && !f[320]; // c2t62i6
	assign leaf[102] = !f[346] && f[543] && f[154] && f[320]; // c2t62i6
	assign leaf[103] = f[346] && !f[582] && !f[527] && !f[637]; // c2t62i6
	assign leaf[104] = f[346] && !f[582] && !f[527] && f[637]; // c2t62i6
	assign leaf[105] = f[346] && !f[582] && f[527] && !f[604]; // c2t62i6
	assign leaf[106] = f[346] && !f[582] && f[527] && f[604]; // c2t62i6
	assign leaf[107] = f[346] && f[582] && !f[633] && !f[522]; // c2t62i6
	assign leaf[108] = f[346] && f[582] && !f[633] && f[522]; // c2t62i6
	assign leaf[109] = f[346] && f[582] && f[633] && !f[547]; // c2t62i6
	assign leaf[110] = f[346] && f[582] && f[633] && f[547]; // c2t62i6
	assign leaf[111] = !f[319] && !f[344] && !f[321] && !f[127]; // c2t72i7
	assign leaf[112] = !f[319] && !f[344] && !f[321] && f[127]; // c2t72i7
	assign leaf[113] = !f[319] && !f[344] && f[321] && !f[499]; // c2t72i7
	assign leaf[114] = !f[319] && !f[344] && f[321] && f[499]; // c2t72i7
	assign leaf[115] = !f[319] && f[344] && !f[316] && !f[425]; // c2t72i7
	assign leaf[116] = !f[319] && f[344] && !f[316] && f[425]; // c2t72i7
	assign leaf[117] = !f[319] && f[344] && f[316] && !f[372]; // c2t72i7
	assign leaf[118] = !f[319] && f[344] && f[316] && f[372]; // c2t72i7
	assign leaf[119] = f[319] && !f[473] && !f[581] && !f[527]; // c2t72i7
	assign leaf[120] = f[319] && !f[473] && !f[581] && f[527]; // c2t72i7
	assign leaf[121] = f[319] && !f[473] && f[581] && !f[490]; // c2t72i7
	assign leaf[122] = f[319] && !f[473] && f[581] && f[490]; // c2t72i7
	assign leaf[123] = f[319] && f[473] && !f[454] && !f[539]; // c2t72i7
	assign leaf[124] = f[319] && f[473] && !f[454] && f[539]; // c2t72i7
	assign leaf[125] = f[319] && f[473] && f[454]; // c2t72i7
	assign leaf[126] = !f[543] && !f[125] && !f[511] && !f[501]; // c2t82i8
	assign leaf[127] = !f[543] && !f[125] && !f[511] && f[501]; // c2t82i8
	assign leaf[128] = !f[543] && !f[125] && f[511] && !f[630]; // c2t82i8
	assign leaf[129] = !f[543] && !f[125] && f[511] && f[630]; // c2t82i8
	assign leaf[130] = !f[543] && f[125] && !f[458] && !f[631]; // c2t82i8
	assign leaf[131] = !f[543] && f[125] && !f[458] && f[631]; // c2t82i8
	assign leaf[132] = !f[543] && f[125] && f[458] && !f[659]; // c2t82i8
	assign leaf[133] = !f[543] && f[125] && f[458] && f[659]; // c2t82i8
	assign leaf[134] = f[543] && !f[607] && !f[524] && !f[470]; // c2t82i8
	assign leaf[135] = f[543] && !f[607] && !f[524] && f[470]; // c2t82i8
	assign leaf[136] = f[543] && !f[607] && f[524] && !f[344]; // c2t82i8
	assign leaf[137] = f[543] && !f[607] && f[524] && f[344]; // c2t82i8
	assign leaf[138] = f[543] && f[607] && !f[496] && !f[442]; // c2t82i8
	assign leaf[139] = f[543] && f[607] && !f[496] && f[442]; // c2t82i8
	assign leaf[140] = f[543] && f[607] && f[496] && !f[594]; // c2t82i8
	assign leaf[141] = f[543] && f[607] && f[496] && f[594]; // c2t82i8
	assign leaf[142] = !f[345] && !f[320] && !f[343] && !f[379]; // c2t92i9
	assign leaf[143] = !f[345] && !f[320] && !f[343] && f[379]; // c2t92i9
	assign leaf[144] = !f[345] && !f[320] && f[343] && !f[399]; // c2t92i9
	assign leaf[145] = !f[345] && !f[320] && f[343] && f[399]; // c2t92i9
	assign leaf[146] = !f[345] && f[320] && !f[554] && !f[473]; // c2t92i9
	assign leaf[147] = !f[345] && f[320] && !f[554] && f[473]; // c2t92i9
	assign leaf[148] = !f[345] && f[320] && f[554] && !f[660]; // c2t92i9
	assign leaf[149] = !f[345] && f[320] && f[554] && f[660]; // c2t92i9
	assign leaf[150] = f[345] && !f[568] && !f[401] && !f[515]; // c2t92i9
	assign leaf[151] = f[345] && !f[568] && !f[401] && f[515]; // c2t92i9
	assign leaf[152] = f[345] && !f[568] && f[401] && !f[511]; // c2t92i9
	assign leaf[153] = f[345] && !f[568] && f[401] && f[511]; // c2t92i9
	assign leaf[154] = f[345] && f[568] && !f[464] && !f[622]; // c2t92i9
	assign leaf[155] = f[345] && f[568] && !f[464] && f[622]; // c2t92i9
	assign leaf[156] = f[345] && f[568] && f[464] && !f[658]; // c2t92i9
	assign leaf[157] = f[345] && f[568] && f[464] && f[658]; // c2t92i9
	assign leaf[158] = !f[151] && !f[657] && !f[156] && !f[527]; // c2t102i10
	assign leaf[159] = !f[151] && !f[657] && !f[156] && f[527]; // c2t102i10
	assign leaf[160] = !f[151] && !f[657] && f[156] && !f[322]; // c2t102i10
	assign leaf[161] = !f[151] && !f[657] && f[156] && f[322]; // c2t102i10
	assign leaf[162] = !f[151] && f[657] && !f[636] && !f[717]; // c2t102i10
	assign leaf[163] = !f[151] && f[657] && !f[636] && f[717]; // c2t102i10
	assign leaf[164] = !f[151] && f[657] && f[636] && !f[516]; // c2t102i10
	assign leaf[165] = !f[151] && f[657] && f[636] && f[516]; // c2t102i10
	assign leaf[166] = f[151] && !f[317] && !f[545] && !f[487]; // c2t102i10
	assign leaf[167] = f[151] && !f[317] && !f[545] && f[487]; // c2t102i10
	assign leaf[168] = f[151] && !f[317] && f[545] && !f[342]; // c2t102i10
	assign leaf[169] = f[151] && !f[317] && f[545] && f[342]; // c2t102i10
	assign leaf[170] = f[151] && f[317] && !f[639] && !f[372]; // c2t102i10
	assign leaf[171] = f[151] && f[317] && !f[639] && f[372]; // c2t102i10
	assign leaf[172] = f[151] && f[317] && f[639] && !f[554]; // c2t102i10
	assign leaf[173] = f[151] && f[317] && f[639] && f[554]; // c2t102i10
	assign leaf[174] = !f[580] && !f[525] && !f[635] && !f[471]; // c2t112i11
	assign leaf[175] = !f[580] && !f[525] && !f[635] && f[471]; // c2t112i11
	assign leaf[176] = !f[580] && !f[525] && f[635] && !f[551]; // c2t112i11
	assign leaf[177] = !f[580] && !f[525] && f[635] && f[551]; // c2t112i11
	assign leaf[178] = !f[580] && f[525] && !f[605] && !f[387]; // c2t112i11
	assign leaf[179] = !f[580] && f[525] && !f[605] && f[387]; // c2t112i11
	assign leaf[180] = !f[580] && f[525] && f[605] && !f[434]; // c2t112i11
	assign leaf[181] = !f[580] && f[525] && f[605] && f[434]; // c2t112i11
	assign leaf[182] = f[580] && !f[468] && !f[414] && !f[662]; // c2t112i11
	assign leaf[183] = f[580] && !f[468] && !f[414] && f[662]; // c2t112i11
	assign leaf[184] = f[580] && !f[468] && f[414]; // c2t112i11
	assign leaf[185] = f[580] && f[468] && !f[520] && !f[131]; // c2t112i11
	assign leaf[186] = f[580] && f[468] && !f[520] && f[131]; // c2t112i11
	assign leaf[187] = f[580] && f[468] && f[520] && !f[371]; // c2t112i11
	assign leaf[188] = f[580] && f[468] && f[520] && f[371]; // c2t112i11
	assign leaf[189] = !f[128] && !f[149] && !f[516] && !f[473]; // c2t122i12
	assign leaf[190] = !f[128] && !f[149] && !f[516] && f[473]; // c2t122i12
	assign leaf[191] = !f[128] && !f[149] && f[516] && !f[526]; // c2t122i12
	assign leaf[192] = !f[128] && !f[149] && f[516] && f[526]; // c2t122i12
	assign leaf[193] = !f[128] && f[149] && !f[317] && !f[259]; // c2t122i12
	assign leaf[194] = !f[128] && f[149] && !f[317] && f[259]; // c2t122i12
	assign leaf[195] = !f[128] && f[149] && f[317] && !f[155]; // c2t122i12
	assign leaf[196] = !f[128] && f[149] && f[317] && f[155]; // c2t122i12
	assign leaf[197] = f[128] && !f[630] && !f[294] && !f[292]; // c2t122i12
	assign leaf[198] = f[128] && !f[630] && !f[294] && f[292]; // c2t122i12
	assign leaf[199] = f[128] && !f[630] && f[294] && !f[607]; // c2t122i12
	assign leaf[200] = f[128] && !f[630] && f[294] && f[607]; // c2t122i12
	assign leaf[201] = f[128] && f[630] && !f[487] && !f[352]; // c2t122i12
	assign leaf[202] = f[128] && f[630] && !f[487] && f[352]; // c2t122i12
	assign leaf[203] = f[128] && f[630] && f[487] && !f[464]; // c2t122i12
	assign leaf[204] = f[128] && f[630] && f[487] && f[464]; // c2t122i12
	assign leaf[205] = !f[345] && !f[348] && !f[370] && !f[607]; // c2t132i13
	assign leaf[206] = !f[345] && !f[348] && !f[370] && f[607]; // c2t132i13
	assign leaf[207] = !f[345] && !f[348] && f[370] && !f[342]; // c2t132i13
	assign leaf[208] = !f[345] && !f[348] && f[370] && f[342]; // c2t132i13
	assign leaf[209] = !f[345] && f[348] && !f[581] && !f[526]; // c2t132i13
	assign leaf[210] = !f[345] && f[348] && !f[581] && f[526]; // c2t132i13
	assign leaf[211] = !f[345] && f[348] && f[581] && !f[440]; // c2t132i13
	assign leaf[212] = !f[345] && f[348] && f[581] && f[440]; // c2t132i13
	assign leaf[213] = f[345] && !f[401] && !f[515] && !f[186]; // c2t132i13
	assign leaf[214] = f[345] && !f[401] && !f[515] && f[186]; // c2t132i13
	assign leaf[215] = f[345] && !f[401] && f[515] && !f[293]; // c2t132i13
	assign leaf[216] = f[345] && !f[401] && f[515] && f[293]; // c2t132i13
	assign leaf[217] = f[345] && f[401] && !f[317] && !f[292]; // c2t132i13
	assign leaf[218] = f[345] && f[401] && !f[317] && f[292]; // c2t132i13
	assign leaf[219] = f[345] && f[401] && f[317] && !f[667]; // c2t132i13
	assign leaf[220] = f[345] && f[401] && f[317] && f[667]; // c2t132i13
	assign leaf[221] = !f[683] && !f[659] && !f[492] && !f[576]; // c2t142i14
	assign leaf[222] = !f[683] && !f[659] && !f[492] && f[576]; // c2t142i14
	assign leaf[223] = !f[683] && !f[659] && f[492] && !f[352]; // c2t142i14
	assign leaf[224] = !f[683] && !f[659] && f[492] && f[352]; // c2t142i14
	assign leaf[225] = !f[683] && f[659] && !f[544] && !f[514]; // c2t142i14
	assign leaf[226] = !f[683] && f[659] && !f[544] && f[514]; // c2t142i14
	assign leaf[227] = !f[683] && f[659] && f[544] && !f[494]; // c2t142i14
	assign leaf[228] = !f[683] && f[659] && f[544] && f[494]; // c2t142i14
	assign leaf[229] = f[683] && !f[403] && !f[691] && !f[598]; // c2t142i14
	assign leaf[230] = f[683] && !f[403] && !f[691] && f[598]; // c2t142i14
	assign leaf[231] = f[683] && !f[403] && f[691]; // c2t142i14
	assign leaf[232] = f[683] && f[403] && !f[610]; // c2t142i14
	assign leaf[233] = f[683] && f[403] && f[610] && !f[325]; // c2t142i14
	assign leaf[234] = f[683] && f[403] && f[610] && f[325]; // c2t142i14
	assign leaf[235] = !f[345] && !f[348] && !f[342] && !f[455]; // c2t152i15
	assign leaf[236] = !f[345] && !f[348] && !f[342] && f[455]; // c2t152i15
	assign leaf[237] = !f[345] && !f[348] && f[342] && !f[398]; // c2t152i15
	assign leaf[238] = !f[345] && !f[348] && f[342] && f[398]; // c2t152i15
	assign leaf[239] = !f[345] && f[348] && !f[444] && !f[580]; // c2t152i15
	assign leaf[240] = !f[345] && f[348] && !f[444] && f[580]; // c2t152i15
	assign leaf[241] = !f[345] && f[348] && f[444] && !f[386]; // c2t152i15
	assign leaf[242] = !f[345] && f[348] && f[444] && f[386]; // c2t152i15
	assign leaf[243] = f[345] && !f[401] && !f[515] && !f[351]; // c2t152i15
	assign leaf[244] = f[345] && !f[401] && !f[515] && f[351]; // c2t152i15
	assign leaf[245] = f[345] && !f[401] && f[515] && !f[427]; // c2t152i15
	assign leaf[246] = f[345] && !f[401] && f[515] && f[427]; // c2t152i15
	assign leaf[247] = f[345] && f[401] && !f[290] && !f[482]; // c2t152i15
	assign leaf[248] = f[345] && f[401] && !f[290] && f[482]; // c2t152i15
	assign leaf[249] = f[345] && f[401] && f[290] && !f[667]; // c2t152i15
	assign leaf[250] = f[345] && f[401] && f[290] && f[667]; // c2t152i15
	assign leaf[251] = !f[150] && !f[657] && !f[157] && !f[471]; // c2t162i16
	assign leaf[252] = !f[150] && !f[657] && !f[157] && f[471]; // c2t162i16
	assign leaf[253] = !f[150] && !f[657] && f[157] && !f[322]; // c2t162i16
	assign leaf[254] = !f[150] && !f[657] && f[157] && f[322]; // c2t162i16
	assign leaf[255] = !f[150] && f[657] && !f[403] && !f[663]; // c2t162i16
	assign leaf[256] = !f[150] && f[657] && !f[403] && f[663]; // c2t162i16
	assign leaf[257] = !f[150] && f[657] && f[403] && !f[125]; // c2t162i16
	assign leaf[258] = !f[150] && f[657] && f[403] && f[125]; // c2t162i16
	assign leaf[259] = f[150] && !f[290] && !f[315] && !f[409]; // c2t162i16
	assign leaf[260] = f[150] && !f[290] && !f[315] && f[409]; // c2t162i16
	assign leaf[261] = f[150] && !f[290] && f[315] && !f[399]; // c2t162i16
	assign leaf[262] = f[150] && !f[290] && f[315] && f[399]; // c2t162i16
	assign leaf[263] = f[150] && f[290] && !f[269] && !f[538]; // c2t162i16
	assign leaf[264] = f[150] && f[290] && !f[269] && f[538]; // c2t162i16
	assign leaf[265] = f[150] && f[290] && f[269] && !f[625]; // c2t162i16
	assign leaf[266] = f[150] && f[290] && f[269] && f[625]; // c2t162i16
	assign leaf[267] = !f[514] && !f[379] && !f[319] && !f[546]; // c2t172i17
	assign leaf[268] = !f[514] && !f[379] && !f[319] && f[546]; // c2t172i17
	assign leaf[269] = !f[514] && !f[379] && f[319] && !f[570]; // c2t172i17
	assign leaf[270] = !f[514] && !f[379] && f[319] && f[570]; // c2t172i17
	assign leaf[271] = !f[514] && f[379] && !f[516] && !f[454]; // c2t172i17
	assign leaf[272] = !f[514] && f[379] && !f[516] && f[454]; // c2t172i17
	assign leaf[273] = !f[514] && f[379] && f[516] && !f[607]; // c2t172i17
	assign leaf[274] = !f[514] && f[379] && f[516] && f[607]; // c2t172i17
	assign leaf[275] = f[514] && !f[343] && !f[580] && !f[635]; // c2t172i17
	assign leaf[276] = f[514] && !f[343] && !f[580] && f[635]; // c2t172i17
	assign leaf[277] = f[514] && !f[343] && f[580] && !f[468]; // c2t172i17
	assign leaf[278] = f[514] && !f[343] && f[580] && f[468]; // c2t172i17
	assign leaf[279] = f[514] && f[343] && !f[427] && !f[401]; // c2t172i17
	assign leaf[280] = f[514] && f[343] && !f[427] && f[401]; // c2t172i17
	assign leaf[281] = f[514] && f[343] && f[427] && !f[375]; // c2t172i17
	assign leaf[282] = f[514] && f[343] && f[427] && f[375]; // c2t172i17
	assign leaf[283] = !f[513] && !f[377] && !f[572] && !f[509]; // c2t182i18
	assign leaf[284] = !f[513] && !f[377] && !f[572] && f[509]; // c2t182i18
	assign leaf[285] = !f[513] && !f[377] && f[572] && !f[634]; // c2t182i18
	assign leaf[286] = !f[513] && !f[377] && f[572] && f[634]; // c2t182i18
	assign leaf[287] = !f[513] && f[377] && !f[454] && !f[487]; // c2t182i18
	assign leaf[288] = !f[513] && f[377] && !f[454] && f[487]; // c2t182i18
	assign leaf[289] = !f[513] && f[377] && f[454] && !f[492]; // c2t182i18
	assign leaf[290] = !f[513] && f[377] && f[454] && f[492]; // c2t182i18
	assign leaf[291] = f[513] && !f[370] && !f[373] && !f[348]; // c2t182i18
	assign leaf[292] = f[513] && !f[370] && !f[373] && f[348]; // c2t182i18
	assign leaf[293] = f[513] && !f[370] && f[373] && !f[318]; // c2t182i18
	assign leaf[294] = f[513] && !f[370] && f[373] && f[318]; // c2t182i18
	assign leaf[295] = f[513] && f[370] && !f[260] && !f[405]; // c2t182i18
	assign leaf[296] = f[513] && f[370] && !f[260] && f[405]; // c2t182i18
	assign leaf[297] = f[513] && f[370] && f[260] && !f[398]; // c2t182i18
	assign leaf[298] = f[513] && f[370] && f[260] && f[398]; // c2t182i18
	assign leaf[299] = !f[373] && !f[458] && !f[377] && !f[176]; // c2t192i19
	assign leaf[300] = !f[373] && !f[458] && !f[377] && f[176]; // c2t192i19
	assign leaf[301] = !f[373] && !f[458] && f[377] && !f[429]; // c2t192i19
	assign leaf[302] = !f[373] && !f[458] && f[377] && f[429]; // c2t192i19
	assign leaf[303] = !f[373] && f[458] && !f[685] && !f[381]; // c2t192i19
	assign leaf[304] = !f[373] && f[458] && !f[685] && f[381]; // c2t192i19
	assign leaf[305] = !f[373] && f[458] && f[685] && !f[599]; // c2t192i19
	assign leaf[306] = !f[373] && f[458] && f[685] && f[599]; // c2t192i19
	assign leaf[307] = f[373] && !f[453] && !f[97] && !f[501]; // c2t192i19
	assign leaf[308] = f[373] && !f[453] && !f[97] && f[501]; // c2t192i19
	assign leaf[309] = f[373] && !f[453] && f[97] && !f[290]; // c2t192i19
	assign leaf[310] = f[373] && !f[453] && f[97] && f[290]; // c2t192i19
	assign leaf[311] = f[373] && f[453] && !f[291] && !f[295]; // c2t192i19
	assign leaf[312] = f[373] && f[453] && !f[291] && f[295]; // c2t192i19
	assign leaf[313] = f[373] && f[453] && f[291] && !f[581]; // c2t192i19
	assign leaf[314] = f[373] && f[453] && f[291] && f[581]; // c2t192i19
	assign leaf[315] = !f[682] && !f[488] && !f[380] && !f[547]; // c2t202i20
	assign leaf[316] = !f[682] && !f[488] && !f[380] && f[547]; // c2t202i20
	assign leaf[317] = !f[682] && !f[488] && f[380] && !f[517]; // c2t202i20
	assign leaf[318] = !f[682] && !f[488] && f[380] && f[517]; // c2t202i20
	assign leaf[319] = !f[682] && f[488] && !f[389] && !f[508]; // c2t202i20
	assign leaf[320] = !f[682] && f[488] && !f[389] && f[508]; // c2t202i20
	assign leaf[321] = !f[682] && f[488] && f[389] && !f[269]; // c2t202i20
	assign leaf[322] = !f[682] && f[488] && f[389] && f[269]; // c2t202i20
	assign leaf[323] = f[682] && !f[658] && !f[577] && !f[387]; // c2t202i20
	assign leaf[324] = f[682] && !f[658] && !f[577] && f[387]; // c2t202i20
	assign leaf[325] = f[682] && !f[658] && f[577] && !f[545]; // c2t202i20
	assign leaf[326] = f[682] && !f[658] && f[577] && f[545]; // c2t202i20
	assign leaf[327] = f[682] && f[658] && !f[404] && !f[570]; // c2t202i20
	assign leaf[328] = f[682] && f[658] && !f[404] && f[570]; // c2t202i20
	assign leaf[329] = f[682] && f[658] && f[404] && !f[541]; // c2t202i20
	assign leaf[330] = f[682] && f[658] && f[404] && f[541]; // c2t202i20
	assign leaf[331] = !f[152] && !f[417] && !f[98] && !f[500]; // c2t212i21
	assign leaf[332] = !f[152] && !f[417] && !f[98] && f[500]; // c2t212i21
	assign leaf[333] = !f[152] && !f[417] && f[98] && !f[292]; // c2t212i21
	assign leaf[334] = !f[152] && !f[417] && f[98] && f[292]; // c2t212i21
	assign leaf[335] = !f[152] && f[417] && !f[343] && !f[240]; // c2t212i21
	assign leaf[336] = !f[152] && f[417] && !f[343] && f[240]; // c2t212i21
	assign leaf[337] = !f[152] && f[417] && f[343]; // c2t212i21
	assign leaf[338] = f[152] && !f[291] && !f[315] && !f[637]; // c2t212i21
	assign leaf[339] = f[152] && !f[291] && !f[315] && f[637]; // c2t212i21
	assign leaf[340] = f[152] && !f[291] && f[315] && !f[655]; // c2t212i21
	assign leaf[341] = f[152] && !f[291] && f[315] && f[655]; // c2t212i21
	assign leaf[342] = f[152] && f[291] && !f[547] && !f[462]; // c2t212i21
	assign leaf[343] = f[152] && f[291] && !f[547] && f[462]; // c2t212i21
	assign leaf[344] = f[152] && f[291] && f[547] && !f[240]; // c2t212i21
	assign leaf[345] = f[152] && f[291] && f[547] && f[240]; // c2t212i21
	assign leaf[346] = !f[380] && !f[397] && !f[372] && !f[204]; // c2t222i22
	assign leaf[347] = !f[380] && !f[397] && !f[372] && f[204]; // c2t222i22
	assign leaf[348] = !f[380] && !f[397] && f[372] && !f[377]; // c2t222i22
	assign leaf[349] = !f[380] && !f[397] && f[372] && f[377]; // c2t222i22
	assign leaf[350] = !f[380] && f[397] && !f[405] && !f[451]; // c2t222i22
	assign leaf[351] = !f[380] && f[397] && !f[405] && f[451]; // c2t222i22
	assign leaf[352] = !f[380] && f[397] && f[405] && !f[159]; // c2t222i22
	assign leaf[353] = !f[380] && f[397] && f[405] && f[159]; // c2t222i22
	assign leaf[354] = f[380] && !f[438] && !f[634] && !f[579]; // c2t222i22
	assign leaf[355] = f[380] && !f[438] && !f[634] && f[579]; // c2t222i22
	assign leaf[356] = f[380] && !f[438] && f[634] && !f[493]; // c2t222i22
	assign leaf[357] = f[380] && !f[438] && f[634] && f[493]; // c2t222i22
	assign leaf[358] = f[380] && f[438] && !f[511] && !f[499]; // c2t222i22
	assign leaf[359] = f[380] && f[438] && !f[511] && f[499]; // c2t222i22
	assign leaf[360] = f[380] && f[438] && f[511] && !f[630]; // c2t222i22
	assign leaf[361] = f[380] && f[438] && f[511] && f[630]; // c2t222i22
	assign leaf[362] = !f[685] && !f[353] && !f[122] && !f[566]; // c2t232i23
	assign leaf[363] = !f[685] && !f[353] && !f[122] && f[566]; // c2t232i23
	assign leaf[364] = !f[685] && !f[353] && f[122] && !f[318]; // c2t232i23
	assign leaf[365] = !f[685] && !f[353] && f[122] && f[318]; // c2t232i23
	assign leaf[366] = !f[685] && f[353] && !f[322] && !f[356]; // c2t232i23
	assign leaf[367] = !f[685] && f[353] && !f[322] && f[356]; // c2t232i23
	assign leaf[368] = !f[685] && f[353] && f[322] && !f[582]; // c2t232i23
	assign leaf[369] = !f[685] && f[353] && f[322] && f[582]; // c2t232i23
	assign leaf[370] = f[685] && !f[665] && !f[717] && !f[376]; // c2t232i23
	assign leaf[371] = f[685] && !f[665] && !f[717] && f[376]; // c2t232i23
	assign leaf[372] = f[685] && !f[665] && f[717]; // c2t232i23
	assign leaf[373] = f[685] && f[665] && !f[582] && !f[463]; // c2t232i23
	assign leaf[374] = f[685] && f[665] && !f[582] && f[463]; // c2t232i23
	assign leaf[375] = f[685] && f[665] && f[582]; // c2t232i23
	assign leaf[376] = !f[501] && !f[373] && !f[349] && !f[398]; // c2t242i24
	assign leaf[377] = !f[501] && !f[373] && !f[349] && f[398]; // c2t242i24
	assign leaf[378] = !f[501] && !f[373] && f[349] && !f[415]; // c2t242i24
	assign leaf[379] = !f[501] && !f[373] && f[349] && f[415]; // c2t242i24
	assign leaf[380] = !f[501] && f[373] && !f[426] && !f[547]; // c2t242i24
	assign leaf[381] = !f[501] && f[373] && !f[426] && f[547]; // c2t242i24
	assign leaf[382] = !f[501] && f[373] && f[426] && !f[290]; // c2t242i24
	assign leaf[383] = !f[501] && f[373] && f[426] && f[290]; // c2t242i24
	assign leaf[384] = f[501] && !f[370] && !f[654] && !f[264]; // c2t242i24
	assign leaf[385] = f[501] && !f[370] && !f[654] && f[264]; // c2t242i24
	assign leaf[386] = f[501] && !f[370] && f[654]; // c2t242i24
	assign leaf[387] = f[501] && f[370]; // c2t242i24
	assign leaf[388] = !f[352] && !f[566] && !f[407] && !f[371]; // c2t252i25
	assign leaf[389] = !f[352] && !f[566] && !f[407] && f[371]; // c2t252i25
	assign leaf[390] = !f[352] && !f[566] && f[407] && !f[512]; // c2t252i25
	assign leaf[391] = !f[352] && !f[566] && f[407] && f[512]; // c2t252i25
	assign leaf[392] = !f[352] && f[566] && !f[342] && !f[301]; // c2t252i25
	assign leaf[393] = !f[352] && f[566] && !f[342] && f[301]; // c2t252i25
	assign leaf[394] = !f[352] && f[566] && f[342] && !f[298]; // c2t252i25
	assign leaf[395] = !f[352] && f[566] && f[342] && f[298]; // c2t252i25
	assign leaf[396] = f[352] && !f[411] && !f[579] && !f[635]; // c2t252i25
	assign leaf[397] = f[352] && !f[411] && !f[579] && f[635]; // c2t252i25
	assign leaf[398] = f[352] && !f[411] && f[579] && !f[466]; // c2t252i25
	assign leaf[399] = f[352] && !f[411] && f[579] && f[466]; // c2t252i25
	assign leaf[400] = f[352] && f[411] && !f[388] && !f[445]; // c2t252i25
	assign leaf[401] = f[352] && f[411] && !f[388] && f[445]; // c2t252i25
	assign leaf[402] = f[352] && f[411] && f[388] && !f[234]; // c2t252i25
	assign leaf[403] = f[352] && f[411] && f[388] && f[234]; // c2t252i25
	assign leaf[404] = !f[152] && !f[497] && !f[580] && !f[415]; // c2t262i26
	assign leaf[405] = !f[152] && !f[497] && !f[580] && f[415]; // c2t262i26
	assign leaf[406] = !f[152] && !f[497] && f[580] && !f[260]; // c2t262i26
	assign leaf[407] = !f[152] && !f[497] && f[580] && f[260]; // c2t262i26
	assign leaf[408] = !f[152] && f[497] && !f[605] && !f[636]; // c2t262i26
	assign leaf[409] = !f[152] && f[497] && !f[605] && f[636]; // c2t262i26
	assign leaf[410] = !f[152] && f[497] && f[605] && !f[437]; // c2t262i26
	assign leaf[411] = !f[152] && f[497] && f[605] && f[437]; // c2t262i26
	assign leaf[412] = f[152] && !f[409] && !f[464] && !f[355]; // c2t262i26
	assign leaf[413] = f[152] && !f[409] && !f[464] && f[355]; // c2t262i26
	assign leaf[414] = f[152] && !f[409] && f[464] && !f[440]; // c2t262i26
	assign leaf[415] = f[152] && !f[409] && f[464] && f[440]; // c2t262i26
	assign leaf[416] = f[152] && f[409] && !f[519] && !f[438]; // c2t262i26
	assign leaf[417] = f[152] && f[409] && !f[519] && f[438]; // c2t262i26
	assign leaf[418] = f[152] && f[409] && f[519] && !f[609]; // c2t262i26
	assign leaf[419] = f[152] && f[409] && f[519] && f[609]; // c2t262i26
	assign leaf[420] = !f[372] && !f[347] && !f[397] && !f[679]; // c2t272i27
	assign leaf[421] = !f[372] && !f[347] && !f[397] && f[679]; // c2t272i27
	assign leaf[422] = !f[372] && !f[347] && f[397] && !f[313]; // c2t272i27
	assign leaf[423] = !f[372] && !f[347] && f[397] && f[313]; // c2t272i27
	assign leaf[424] = !f[372] && f[347] && !f[444] && !f[580]; // c2t272i27
	assign leaf[425] = !f[372] && f[347] && !f[444] && f[580]; // c2t272i27
	assign leaf[426] = !f[372] && f[347] && f[444] && !f[567]; // c2t272i27
	assign leaf[427] = !f[372] && f[347] && f[444] && f[567]; // c2t272i27
	assign leaf[428] = f[372] && !f[316] && !f[291] && !f[482]; // c2t272i27
	assign leaf[429] = f[372] && !f[316] && !f[291] && f[482]; // c2t272i27
	assign leaf[430] = f[372] && !f[316] && f[291] && !f[444]; // c2t272i27
	assign leaf[431] = f[372] && !f[316] && f[291] && f[444]; // c2t272i27
	assign leaf[432] = f[372] && f[316] && !f[400] && !f[515]; // c2t272i27
	assign leaf[433] = f[372] && f[316] && !f[400] && f[515]; // c2t272i27
	assign leaf[434] = f[372] && f[316] && f[400] && !f[652]; // c2t272i27
	assign leaf[435] = f[372] && f[316] && f[400] && f[652]; // c2t272i27
	assign leaf[436] = !f[514] && !f[379] && !f[572] && !f[174]; // c2t282i28
	assign leaf[437] = !f[514] && !f[379] && !f[572] && f[174]; // c2t282i28
	assign leaf[438] = !f[514] && !f[379] && f[572] && !f[294]; // c2t282i28
	assign leaf[439] = !f[514] && !f[379] && f[572] && f[294]; // c2t282i28
	assign leaf[440] = !f[514] && f[379] && !f[517] && !f[427]; // c2t282i28
	assign leaf[441] = !f[514] && f[379] && !f[517] && f[427]; // c2t282i28
	assign leaf[442] = !f[514] && f[379] && f[517] && !f[215]; // c2t282i28
	assign leaf[443] = !f[514] && f[379] && f[517] && f[215]; // c2t282i28
	assign leaf[444] = f[514] && !f[460] && !f[624] && !f[404]; // c2t282i28
	assign leaf[445] = f[514] && !f[460] && !f[624] && f[404]; // c2t282i28
	assign leaf[446] = f[514] && !f[460] && f[624] && !f[545]; // c2t282i28
	assign leaf[447] = f[514] && !f[460] && f[624] && f[545]; // c2t282i28
	assign leaf[448] = f[514] && f[460] && !f[679] && !f[409]; // c2t282i28
	assign leaf[449] = f[514] && f[460] && !f[679] && f[409]; // c2t282i28
	assign leaf[450] = f[514] && f[460] && f[679] && !f[631]; // c2t282i28
	assign leaf[451] = f[514] && f[460] && f[679] && f[631]; // c2t282i28
	assign leaf[452] = !f[473] && !f[514] && !f[379] && !f[548]; // c2t292i29
	assign leaf[453] = !f[473] && !f[514] && !f[379] && f[548]; // c2t292i29
	assign leaf[454] = !f[473] && !f[514] && f[379] && !f[638]; // c2t292i29
	assign leaf[455] = !f[473] && !f[514] && f[379] && f[638]; // c2t292i29
	assign leaf[456] = !f[473] && f[514] && !f[433] && !f[353]; // c2t292i29
	assign leaf[457] = !f[473] && f[514] && !f[433] && f[353]; // c2t292i29
	assign leaf[458] = !f[473] && f[514] && f[433] && !f[651]; // c2t292i29
	assign leaf[459] = !f[473] && f[514] && f[433] && f[651]; // c2t292i29
	assign leaf[460] = f[473] && !f[343] && !f[354]; // c2t292i29
	assign leaf[461] = f[473] && !f[343] && f[354]; // c2t292i29
	assign leaf[462] = f[473] && f[343]; // c2t292i29
	assign leaf[463] = !f[682] && !f[713] && !f[372] && !f[351]; // c2t302i30
	assign leaf[464] = !f[682] && !f[713] && !f[372] && f[351]; // c2t302i30
	assign leaf[465] = !f[682] && !f[713] && f[372] && !f[316]; // c2t302i30
	assign leaf[466] = !f[682] && !f[713] && f[372] && f[316]; // c2t302i30
	assign leaf[467] = !f[682] && f[713] && !f[599]; // c2t302i30
	assign leaf[468] = !f[682] && f[713] && f[599]; // c2t302i30
	assign leaf[469] = f[682] && !f[180] && !f[605]; // c2t302i30
	assign leaf[470] = f[682] && !f[180] && f[605]; // c2t302i30
	assign leaf[471] = f[682] && f[180] && !f[431] && !f[406]; // c2t302i30
	assign leaf[472] = f[682] && f[180] && !f[431] && f[406]; // c2t302i30
	assign leaf[473] = f[682] && f[180] && f[431] && !f[541]; // c2t302i30
	assign leaf[474] = f[682] && f[180] && f[431] && f[541]; // c2t302i30
	assign leaf[475] = !f[176] && !f[485] && !f[516] && !f[455]; // c2t312i31
	assign leaf[476] = !f[176] && !f[485] && !f[516] && f[455]; // c2t312i31
	assign leaf[477] = !f[176] && !f[485] && f[516] && !f[609]; // c2t312i31
	assign leaf[478] = !f[176] && !f[485] && f[516] && f[609]; // c2t312i31
	assign leaf[479] = !f[176] && f[485] && !f[432] && !f[595]; // c2t312i31
	assign leaf[480] = !f[176] && f[485] && !f[432] && f[595]; // c2t312i31
	assign leaf[481] = !f[176] && f[485] && f[432] && !f[685]; // c2t312i31
	assign leaf[482] = !f[176] && f[485] && f[432] && f[685]; // c2t312i31
	assign leaf[483] = f[176] && !f[551] && !f[691] && !f[341]; // c2t312i31
	assign leaf[484] = f[176] && !f[551] && !f[691] && f[341]; // c2t312i31
	assign leaf[485] = f[176] && !f[551] && f[691] && !f[610]; // c2t312i31
	assign leaf[486] = f[176] && !f[551] && f[691] && f[610]; // c2t312i31
	assign leaf[487] = f[176] && f[551] && !f[661] && !f[208]; // c2t312i31
	assign leaf[488] = f[176] && f[551] && !f[661] && f[208]; // c2t312i31
	assign leaf[489] = f[176] && f[551] && f[661] && !f[380]; // c2t312i31
	assign leaf[490] = f[176] && f[551] && f[661] && f[380]; // c2t312i31
	assign leaf[491] = !f[121] && !f[545] && !f[509] && !f[417]; // c2t322i32
	assign leaf[492] = !f[121] && !f[545] && !f[509] && f[417]; // c2t322i32
	assign leaf[493] = !f[121] && !f[545] && f[509] && !f[434]; // c2t322i32
	assign leaf[494] = !f[121] && !f[545] && f[509] && f[434]; // c2t322i32
	assign leaf[495] = !f[121] && f[545] && !f[634] && !f[551]; // c2t322i32
	assign leaf[496] = !f[121] && f[545] && !f[634] && f[551]; // c2t322i32
	assign leaf[497] = !f[121] && f[545] && f[634] && !f[495]; // c2t322i32
	assign leaf[498] = !f[121] && f[545] && f[634] && f[495]; // c2t322i32
	assign leaf[499] = f[121] && !f[232] && !f[290] && !f[605]; // c2t322i32
	assign leaf[500] = f[121] && !f[232] && !f[290] && f[605]; // c2t322i32
	assign leaf[501] = f[121] && !f[232] && f[290]; // c2t322i32
	assign leaf[502] = f[121] && f[232] && !f[496] && !f[181]; // c2t322i32
	assign leaf[503] = f[121] && f[232] && !f[496] && f[181]; // c2t322i32
	assign leaf[504] = f[121] && f[232] && f[496] && !f[633]; // c2t322i32
	assign leaf[505] = f[121] && f[232] && f[496] && f[633]; // c2t322i32
	assign leaf[506] = !f[713] && !f[710] && !f[95] && !f[322]; // c2t332i33
	assign leaf[507] = !f[713] && !f[710] && !f[95] && f[322]; // c2t332i33
	assign leaf[508] = !f[713] && !f[710] && f[95] && !f[262]; // c2t332i33
	assign leaf[509] = !f[713] && !f[710] && f[95] && f[262]; // c2t332i33
	assign leaf[510] = !f[713] && f[710]; // c2t332i33
	assign leaf[511] = f[713] && !f[626]; // c2t332i33
	assign leaf[512] = f[713] && f[626]; // c2t332i33
	assign leaf[513] = !f[639] && !f[677] && !f[351] && !f[372]; // c2t342i34
	assign leaf[514] = !f[639] && !f[677] && !f[351] && f[372]; // c2t342i34
	assign leaf[515] = !f[639] && !f[677] && f[351] && !f[487]; // c2t342i34
	assign leaf[516] = !f[639] && !f[677] && f[351] && f[487]; // c2t342i34
	assign leaf[517] = !f[639] && f[677] && !f[289]; // c2t342i34
	assign leaf[518] = !f[639] && f[677] && f[289]; // c2t342i34
	assign leaf[519] = f[639] && !f[554] && !f[371] && !f[569]; // c2t342i34
	assign leaf[520] = f[639] && !f[554] && !f[371] && f[569]; // c2t342i34
	assign leaf[521] = f[639] && !f[554] && f[371]; // c2t342i34
	assign leaf[522] = f[639] && f[554] && !f[550] && !f[382]; // c2t342i34
	assign leaf[523] = f[639] && f[554] && !f[550] && f[382]; // c2t342i34
	assign leaf[524] = f[639] && f[554] && f[550]; // c2t342i34
	assign leaf[525] = !f[179] && !f[655] && !f[630] && !f[242]; // c2t352i35
	assign leaf[526] = !f[179] && !f[655] && !f[630] && f[242]; // c2t352i35
	assign leaf[527] = !f[179] && !f[655] && f[630] && !f[651]; // c2t352i35
	assign leaf[528] = !f[179] && !f[655] && f[630] && f[651]; // c2t352i35
	assign leaf[529] = !f[179] && f[655] && !f[606] && !f[596]; // c2t352i35
	assign leaf[530] = !f[179] && f[655] && !f[606] && f[596]; // c2t352i35
	assign leaf[531] = !f[179] && f[655] && f[606] && !f[601]; // c2t352i35
	assign leaf[532] = !f[179] && f[655] && f[606] && f[601]; // c2t352i35
	assign leaf[533] = f[179] && !f[599] && !f[341] && !f[666]; // c2t352i35
	assign leaf[534] = f[179] && !f[599] && !f[341] && f[666]; // c2t352i35
	assign leaf[535] = f[179] && !f[599] && f[341] && !f[583]; // c2t352i35
	assign leaf[536] = f[179] && !f[599] && f[341] && f[583]; // c2t352i35
	assign leaf[537] = f[179] && f[599] && !f[690] && !f[409]; // c2t352i35
	assign leaf[538] = f[179] && f[599] && !f[690] && f[409]; // c2t352i35
	assign leaf[539] = f[179] && f[599] && f[690] && !f[636]; // c2t352i35
	assign leaf[540] = f[179] && f[599] && f[690] && f[636]; // c2t352i35
	assign leaf[541] = !f[397] && !f[388] && !f[374] && !f[349]; // c2t362i36
	assign leaf[542] = !f[397] && !f[388] && !f[374] && f[349]; // c2t362i36
	assign leaf[543] = !f[397] && !f[388] && f[374] && !f[318]; // c2t362i36
	assign leaf[544] = !f[397] && !f[388] && f[374] && f[318]; // c2t362i36
	assign leaf[545] = !f[397] && f[388] && !f[399] && !f[214]; // c2t362i36
	assign leaf[546] = !f[397] && f[388] && !f[399] && f[214]; // c2t362i36
	assign leaf[547] = !f[397] && f[388] && f[399] && !f[343]; // c2t362i36
	assign leaf[548] = !f[397] && f[388] && f[399] && f[343]; // c2t362i36
	assign leaf[549] = f[397] && !f[374] && !f[426] && !f[495]; // c2t362i36
	assign leaf[550] = f[397] && !f[374] && !f[426] && f[495]; // c2t362i36
	assign leaf[551] = f[397] && !f[374] && f[426] && !f[508]; // c2t362i36
	assign leaf[552] = f[397] && !f[374] && f[426] && f[508]; // c2t362i36
	assign leaf[553] = f[397] && f[374] && !f[287] && !f[521]; // c2t362i36
	assign leaf[554] = f[397] && f[374] && !f[287] && f[521]; // c2t362i36
	assign leaf[555] = f[397] && f[374] && f[287]; // c2t362i36
	assign leaf[556] = !f[473] && !f[293] && !f[289] && !f[427]; // c2t372i37
	assign leaf[557] = !f[473] && !f[293] && !f[289] && f[427]; // c2t372i37
	assign leaf[558] = !f[473] && !f[293] && f[289] && !f[373]; // c2t372i37
	assign leaf[559] = !f[473] && !f[293] && f[289] && f[373]; // c2t372i37
	assign leaf[560] = !f[473] && f[293] && !f[388] && !f[620]; // c2t372i37
	assign leaf[561] = !f[473] && f[293] && !f[388] && f[620]; // c2t372i37
	assign leaf[562] = !f[473] && f[293] && f[388] && !f[359]; // c2t372i37
	assign leaf[563] = !f[473] && f[293] && f[388] && f[359]; // c2t372i37
	assign leaf[564] = f[473] && !f[416] && !f[485]; // c2t372i37
	assign leaf[565] = f[473] && !f[416] && f[485] && !f[400]; // c2t372i37
	assign leaf[566] = f[473] && !f[416] && f[485] && f[400]; // c2t372i37
	assign leaf[567] = f[473] && f[416]; // c2t372i37
	assign leaf[568] = !f[324] && !f[485] && !f[298] && !f[380]; // c2t382i38
	assign leaf[569] = !f[324] && !f[485] && !f[298] && f[380]; // c2t382i38
	assign leaf[570] = !f[324] && !f[485] && f[298] && !f[432]; // c2t382i38
	assign leaf[571] = !f[324] && !f[485] && f[298] && f[432]; // c2t382i38
	assign leaf[572] = !f[324] && f[485] && !f[285] && !f[343]; // c2t382i38
	assign leaf[573] = !f[324] && f[485] && !f[285] && f[343]; // c2t382i38
	assign leaf[574] = !f[324] && f[485] && f[285] && !f[231]; // c2t382i38
	assign leaf[575] = !f[324] && f[485] && f[285] && f[231]; // c2t382i38
	assign leaf[576] = f[324] && !f[411] && !f[271] && !f[159]; // c2t382i38
	assign leaf[577] = f[324] && !f[411] && !f[271] && f[159]; // c2t382i38
	assign leaf[578] = f[324] && !f[411] && f[271] && !f[606]; // c2t382i38
	assign leaf[579] = f[324] && !f[411] && f[271] && f[606]; // c2t382i38
	assign leaf[580] = f[324] && f[411] && !f[415] && !f[172]; // c2t382i38
	assign leaf[581] = f[324] && f[411] && !f[415] && f[172]; // c2t382i38
	assign leaf[582] = f[324] && f[411] && f[415] && !f[243]; // c2t382i38
	assign leaf[583] = f[324] && f[411] && f[415] && f[243]; // c2t382i38
	assign leaf[584] = !f[95] && !f[547] && !f[630] && !f[652]; // c2t392i39
	assign leaf[585] = !f[95] && !f[547] && !f[630] && f[652]; // c2t392i39
	assign leaf[586] = !f[95] && !f[547] && f[630] && !f[522]; // c2t392i39
	assign leaf[587] = !f[95] && !f[547] && f[630] && f[522]; // c2t392i39
	assign leaf[588] = !f[95] && f[547] && !f[685] && !f[687]; // c2t392i39
	assign leaf[589] = !f[95] && f[547] && !f[685] && f[687]; // c2t392i39
	assign leaf[590] = !f[95] && f[547] && f[685] && !f[461]; // c2t392i39
	assign leaf[591] = !f[95] && f[547] && f[685] && f[461]; // c2t392i39
	assign leaf[592] = f[95] && !f[354] && !f[458] && !f[461]; // c2t392i39
	assign leaf[593] = f[95] && !f[354] && !f[458] && f[461]; // c2t392i39
	assign leaf[594] = f[95] && !f[354] && f[458] && !f[517]; // c2t392i39
	assign leaf[595] = f[95] && !f[354] && f[458] && f[517]; // c2t392i39
	assign leaf[596] = f[95] && f[354] && !f[521]; // c2t392i39
	assign leaf[597] = f[95] && f[354] && f[521] && !f[270]; // c2t392i39
	assign leaf[598] = f[95] && f[354] && f[521] && f[270]; // c2t392i39
	assign leaf[599] = !f[666] && !f[611] && !f[556] && !f[472]; // c2t402i40
	assign leaf[600] = !f[666] && !f[611] && !f[556] && f[472]; // c2t402i40
	assign leaf[601] = !f[666] && !f[611] && f[556] && !f[127]; // c2t402i40
	assign leaf[602] = !f[666] && !f[611] && f[556] && f[127]; // c2t402i40
	assign leaf[603] = !f[666] && f[611] && !f[527] && !f[344]; // c2t402i40
	assign leaf[604] = !f[666] && f[611] && !f[527] && f[344]; // c2t402i40
	assign leaf[605] = !f[666] && f[611] && f[527] && !f[293]; // c2t402i40
	assign leaf[606] = !f[666] && f[611] && f[527] && f[293]; // c2t402i40
	assign leaf[607] = f[666] && !f[525] && !f[582] && !f[576]; // c2t402i40
	assign leaf[608] = f[666] && !f[525] && !f[582] && f[576]; // c2t402i40
	assign leaf[609] = f[666] && !f[525] && f[582]; // c2t402i40
	assign leaf[610] = f[666] && f[525] && !f[155]; // c2t402i40
	assign leaf[611] = f[666] && f[525] && f[155]; // c2t402i40
	assign leaf[612] = !f[409] && !f[354] && !f[97] && !f[149]; // c2t412i41
	assign leaf[613] = !f[409] && !f[354] && !f[97] && f[149]; // c2t412i41
	assign leaf[614] = !f[409] && !f[354] && f[97] && !f[463]; // c2t412i41
	assign leaf[615] = !f[409] && !f[354] && f[97] && f[463]; // c2t412i41
	assign leaf[616] = !f[409] && f[354] && !f[294] && !f[210]; // c2t412i41
	assign leaf[617] = !f[409] && f[354] && !f[294] && f[210]; // c2t412i41
	assign leaf[618] = !f[409] && f[354] && f[294] && !f[371]; // c2t412i41
	assign leaf[619] = !f[409] && f[354] && f[294] && f[371]; // c2t412i41
	assign leaf[620] = f[409] && !f[463] && !f[355] && !f[379]; // c2t412i41
	assign leaf[621] = f[409] && !f[463] && !f[355] && f[379]; // c2t412i41
	assign leaf[622] = f[409] && !f[463] && f[355] && !f[655]; // c2t412i41
	assign leaf[623] = f[409] && !f[463] && f[355] && f[655]; // c2t412i41
	assign leaf[624] = f[409] && f[463] && !f[538] && !f[460]; // c2t412i41
	assign leaf[625] = f[409] && f[463] && !f[538] && f[460]; // c2t412i41
	assign leaf[626] = f[409] && f[463] && f[538] && !f[600]; // c2t412i41
	assign leaf[627] = f[409] && f[463] && f[538] && f[600]; // c2t412i41
	assign leaf[628] = !f[409] && !f[549] && !f[605] && !f[443]; // c2t422i42
	assign leaf[629] = !f[409] && !f[549] && !f[605] && f[443]; // c2t422i42
	assign leaf[630] = !f[409] && !f[549] && f[605] && !f[523]; // c2t422i42
	assign leaf[631] = !f[409] && !f[549] && f[605] && f[523]; // c2t422i42
	assign leaf[632] = !f[409] && f[549] && !f[660] && !f[460]; // c2t422i42
	assign leaf[633] = !f[409] && f[549] && !f[660] && f[460]; // c2t422i42
	assign leaf[634] = !f[409] && f[549] && f[660] && !f[384]; // c2t422i42
	assign leaf[635] = !f[409] && f[549] && f[660] && f[384]; // c2t422i42
	assign leaf[636] = f[409] && !f[463] && !f[176] && !f[681]; // c2t422i42
	assign leaf[637] = f[409] && !f[463] && !f[176] && f[681]; // c2t422i42
	assign leaf[638] = f[409] && !f[463] && f[176] && !f[521]; // c2t422i42
	assign leaf[639] = f[409] && !f[463] && f[176] && f[521]; // c2t422i42
	assign leaf[640] = f[409] && f[463] && !f[609] && !f[201]; // c2t422i42
	assign leaf[641] = f[409] && f[463] && !f[609] && f[201]; // c2t422i42
	assign leaf[642] = f[409] && f[463] && f[609] && !f[469]; // c2t422i42
	assign leaf[643] = f[409] && f[463] && f[609] && f[469]; // c2t422i42
	assign leaf[644] = !f[486] && !f[432] && !f[512] && !f[689]; // c2t432i43
	assign leaf[645] = !f[486] && !f[432] && !f[512] && f[689]; // c2t432i43
	assign leaf[646] = !f[486] && !f[432] && f[512] && !f[404]; // c2t432i43
	assign leaf[647] = !f[486] && !f[432] && f[512] && f[404]; // c2t432i43
	assign leaf[648] = !f[486] && f[432] && !f[455] && !f[403]; // c2t432i43
	assign leaf[649] = !f[486] && f[432] && !f[455] && f[403]; // c2t432i43
	assign leaf[650] = !f[486] && f[432] && f[455] && !f[465]; // c2t432i43
	assign leaf[651] = !f[486] && f[432] && f[455] && f[465]; // c2t432i43
	assign leaf[652] = f[486] && !f[690] && !f[687] && !f[383]; // c2t432i43
	assign leaf[653] = f[486] && !f[690] && !f[687] && f[383]; // c2t432i43
	assign leaf[654] = f[486] && !f[690] && f[687] && !f[598]; // c2t432i43
	assign leaf[655] = f[486] && !f[690] && f[687] && f[598]; // c2t432i43
	assign leaf[656] = f[486] && f[690] && !f[657] && !f[573]; // c2t432i43
	assign leaf[657] = f[486] && f[690] && !f[657] && f[573]; // c2t432i43
	assign leaf[658] = f[486] && f[690] && f[657]; // c2t432i43
	assign leaf[659] = !f[677] && !f[323] && !f[261] && !f[292]; // c2t442i44
	assign leaf[660] = !f[677] && !f[323] && !f[261] && f[292]; // c2t442i44
	assign leaf[661] = !f[677] && !f[323] && f[261] && !f[652]; // c2t442i44
	assign leaf[662] = !f[677] && !f[323] && f[261] && f[652]; // c2t442i44
	assign leaf[663] = !f[677] && f[323] && !f[326] && !f[516]; // c2t442i44
	assign leaf[664] = !f[677] && f[323] && !f[326] && f[516]; // c2t442i44
	assign leaf[665] = !f[677] && f[323] && f[326] && !f[578]; // c2t442i44
	assign leaf[666] = !f[677] && f[323] && f[326] && f[578]; // c2t442i44
	assign leaf[667] = f[677] && !f[158]; // c2t442i44
	assign leaf[668] = f[677] && f[158]; // c2t442i44
	assign leaf[669] = !f[681] && !f[461] && !f[573] && !f[430]; // c2t452i45
	assign leaf[670] = !f[681] && !f[461] && !f[573] && f[430]; // c2t452i45
	assign leaf[671] = !f[681] && !f[461] && f[573] && !f[204]; // c2t452i45
	assign leaf[672] = !f[681] && !f[461] && f[573] && f[204]; // c2t452i45
	assign leaf[673] = !f[681] && f[461] && !f[525] && !f[388]; // c2t452i45
	assign leaf[674] = !f[681] && f[461] && !f[525] && f[388]; // c2t452i45
	assign leaf[675] = !f[681] && f[461] && f[525] && !f[607]; // c2t452i45
	assign leaf[676] = !f[681] && f[461] && f[525] && f[607]; // c2t452i45
	assign leaf[677] = f[681] && !f[603] && !f[686] && !f[462]; // c2t452i45
	assign leaf[678] = f[681] && !f[603] && !f[686] && f[462]; // c2t452i45
	assign leaf[679] = f[681] && !f[603] && f[686] && !f[631]; // c2t452i45
	assign leaf[680] = f[681] && !f[603] && f[686] && f[631]; // c2t452i45
	assign leaf[681] = f[681] && f[603] && !f[432] && !f[685]; // c2t452i45
	assign leaf[682] = f[681] && f[603] && !f[432] && f[685]; // c2t452i45
	assign leaf[683] = f[681] && f[603] && f[432] && !f[594]; // c2t452i45
	assign leaf[684] = f[681] && f[603] && f[432] && f[594]; // c2t452i45
	assign leaf[685] = !f[324] && !f[509] && !f[571] && !f[267]; // c2t462i46
	assign leaf[686] = !f[324] && !f[509] && !f[571] && f[267]; // c2t462i46
	assign leaf[687] = !f[324] && !f[509] && f[571] && !f[297]; // c2t462i46
	assign leaf[688] = !f[324] && !f[509] && f[571] && f[297]; // c2t462i46
	assign leaf[689] = !f[324] && f[509] && !f[457] && !f[403]; // c2t462i46
	assign leaf[690] = !f[324] && f[509] && !f[457] && f[403]; // c2t462i46
	assign leaf[691] = !f[324] && f[509] && f[457] && !f[376]; // c2t462i46
	assign leaf[692] = !f[324] && f[509] && f[457] && f[376]; // c2t462i46
	assign leaf[693] = f[324] && !f[347] && !f[356] && !f[215]; // c2t462i46
	assign leaf[694] = f[324] && !f[347] && !f[356] && f[215]; // c2t462i46
	assign leaf[695] = f[324] && !f[347] && f[356] && !f[204]; // c2t462i46
	assign leaf[696] = f[324] && !f[347] && f[356] && f[204]; // c2t462i46
	assign leaf[697] = f[324] && f[347] && !f[96] && !f[453]; // c2t462i46
	assign leaf[698] = f[324] && f[347] && !f[96] && f[453]; // c2t462i46
	assign leaf[699] = f[324] && f[347] && f[96]; // c2t462i46
	assign leaf[700] = !f[367] && !f[665] && !f[219] && !f[104]; // c2t472i47
	assign leaf[701] = !f[367] && !f[665] && !f[219] && f[104]; // c2t472i47
	assign leaf[702] = !f[367] && !f[665] && f[219] && !f[159]; // c2t472i47
	assign leaf[703] = !f[367] && !f[665] && f[219] && f[159]; // c2t472i47
	assign leaf[704] = !f[367] && f[665] && !f[553] && !f[551]; // c2t472i47
	assign leaf[705] = !f[367] && f[665] && !f[553] && f[551]; // c2t472i47
	assign leaf[706] = !f[367] && f[665] && f[553] && !f[546]; // c2t472i47
	assign leaf[707] = !f[367] && f[665] && f[553] && f[546]; // c2t472i47
	assign leaf[708] = f[367]; // c2t472i47
	assign leaf[709] = !f[418] && !f[473] && !f[571] && !f[510]; // c2t482i48
	assign leaf[710] = !f[418] && !f[473] && !f[571] && f[510]; // c2t482i48
	assign leaf[711] = !f[418] && !f[473] && f[571] && !f[715]; // c2t482i48
	assign leaf[712] = !f[418] && !f[473] && f[571] && f[715]; // c2t482i48
	assign leaf[713] = !f[418] && f[473] && !f[416] && !f[519]; // c2t482i48
	assign leaf[714] = !f[418] && f[473] && !f[416] && f[519]; // c2t482i48
	assign leaf[715] = !f[418] && f[473] && f[416]; // c2t482i48
	assign leaf[716] = f[418]; // c2t482i48
	assign leaf[717] = !f[104] && !f[70] && !f[445] && !f[501]; // c2t492i49
	assign leaf[718] = !f[104] && !f[70] && !f[445] && f[501]; // c2t492i49
	assign leaf[719] = !f[104] && !f[70] && f[445] && !f[552]; // c2t492i49
	assign leaf[720] = !f[104] && !f[70] && f[445] && f[552]; // c2t492i49
	assign leaf[721] = !f[104] && f[70] && !f[152] && !f[493]; // c2t492i49
	assign leaf[722] = !f[104] && f[70] && !f[152] && f[493]; // c2t492i49
	assign leaf[723] = !f[104] && f[70] && f[152]; // c2t492i49
	assign leaf[724] = f[104] && !f[431] && !f[324]; // c2t492i49
	assign leaf[725] = f[104] && !f[431] && f[324]; // c2t492i49
	assign leaf[726] = f[104] && f[431] && !f[322]; // c2t492i49
	assign leaf[727] = f[104] && f[431] && f[322]; // c2t492i49
	assign leaf[728] = !f[95] && !f[390] && !f[235] && !f[351]; // c2t502i50
	assign leaf[729] = !f[95] && !f[390] && !f[235] && f[351]; // c2t502i50
	assign leaf[730] = !f[95] && !f[390] && f[235] && !f[401]; // c2t502i50
	assign leaf[731] = !f[95] && !f[390] && f[235] && f[401]; // c2t502i50
	assign leaf[732] = !f[95] && f[390]; // c2t502i50
	assign leaf[733] = f[95] && !f[262] && !f[453] && !f[402]; // c2t502i50
	assign leaf[734] = f[95] && !f[262] && !f[453] && f[402]; // c2t502i50
	assign leaf[735] = f[95] && !f[262] && f[453]; // c2t502i50
	assign leaf[736] = f[95] && f[262]; // c2t502i50
	assign leaf[737] = !f[134] && !f[411] && !f[356] && !f[470]; // c2t512i51
	assign leaf[738] = !f[134] && !f[411] && !f[356] && f[470]; // c2t512i51
	assign leaf[739] = !f[134] && !f[411] && f[356] && !f[324]; // c2t512i51
	assign leaf[740] = !f[134] && !f[411] && f[356] && f[324]; // c2t512i51
	assign leaf[741] = !f[134] && f[411] && !f[493] && !f[524]; // c2t512i51
	assign leaf[742] = !f[134] && f[411] && !f[493] && f[524]; // c2t512i51
	assign leaf[743] = !f[134] && f[411] && f[493] && !f[515]; // c2t512i51
	assign leaf[744] = !f[134] && f[411] && f[493] && f[515]; // c2t512i51
	assign leaf[745] = f[134] && !f[301]; // c2t512i51
	assign leaf[746] = f[134] && f[301] && !f[467]; // c2t512i51
	assign leaf[747] = f[134] && f[301] && f[467]; // c2t512i51
	assign leaf[748] = !f[708] && !f[514] && !f[432] && !f[231]; // c2t522i52
	assign leaf[749] = !f[708] && !f[514] && !f[432] && f[231]; // c2t522i52
	assign leaf[750] = !f[708] && !f[514] && f[432] && !f[408]; // c2t522i52
	assign leaf[751] = !f[708] && !f[514] && f[432] && f[408]; // c2t522i52
	assign leaf[752] = !f[708] && f[514] && !f[597] && !f[287]; // c2t522i52
	assign leaf[753] = !f[708] && f[514] && !f[597] && f[287]; // c2t522i52
	assign leaf[754] = !f[708] && f[514] && f[597] && !f[184]; // c2t522i52
	assign leaf[755] = !f[708] && f[514] && f[597] && f[184]; // c2t522i52
	assign leaf[756] = f[708] && !f[460]; // c2t522i52
	assign leaf[757] = f[708] && f[460]; // c2t522i52
	assign leaf[758] = !f[242] && !f[154] && !f[213] && !f[299]; // c2t532i53
	assign leaf[759] = !f[242] && !f[154] && !f[213] && f[299]; // c2t532i53
	assign leaf[760] = !f[242] && !f[154] && f[213] && !f[355]; // c2t532i53
	assign leaf[761] = !f[242] && !f[154] && f[213] && f[355]; // c2t532i53
	assign leaf[762] = !f[242] && f[154] && !f[159] && !f[240]; // c2t532i53
	assign leaf[763] = !f[242] && f[154] && !f[159] && f[240]; // c2t532i53
	assign leaf[764] = !f[242] && f[154] && f[159] && !f[358]; // c2t532i53
	assign leaf[765] = !f[242] && f[154] && f[159] && f[358]; // c2t532i53
	assign leaf[766] = f[242] && !f[156] && !f[509] && !f[688]; // c2t532i53
	assign leaf[767] = f[242] && !f[156] && !f[509] && f[688]; // c2t532i53
	assign leaf[768] = f[242] && !f[156] && f[509] && !f[464]; // c2t532i53
	assign leaf[769] = f[242] && !f[156] && f[509] && f[464]; // c2t532i53
	assign leaf[770] = f[242] && f[156] && !f[597] && !f[408]; // c2t532i53
	assign leaf[771] = f[242] && f[156] && !f[597] && f[408]; // c2t532i53
	assign leaf[772] = f[242] && f[156] && f[597] && !f[594]; // c2t532i53
	assign leaf[773] = f[242] && f[156] && f[597] && f[594]; // c2t532i53
	assign leaf[774] = !f[400] && !f[344] && !f[233] && !f[607]; // c2t542i54
	assign leaf[775] = !f[400] && !f[344] && !f[233] && f[607]; // c2t542i54
	assign leaf[776] = !f[400] && !f[344] && f[233] && !f[466]; // c2t542i54
	assign leaf[777] = !f[400] && !f[344] && f[233] && f[466]; // c2t542i54
	assign leaf[778] = !f[400] && f[344] && !f[401] && !f[454]; // c2t542i54
	assign leaf[779] = !f[400] && f[344] && !f[401] && f[454]; // c2t542i54
	assign leaf[780] = !f[400] && f[344] && f[401] && !f[343]; // c2t542i54
	assign leaf[781] = !f[400] && f[344] && f[401] && f[343]; // c2t542i54
	assign leaf[782] = f[400] && !f[376] && !f[372] && !f[432]; // c2t542i54
	assign leaf[783] = f[400] && !f[376] && !f[372] && f[432]; // c2t542i54
	assign leaf[784] = f[400] && !f[376] && f[372] && !f[623]; // c2t542i54
	assign leaf[785] = f[400] && !f[376] && f[372] && f[623]; // c2t542i54
	assign leaf[786] = f[400] && f[376] && !f[659] && !f[295]; // c2t542i54
	assign leaf[787] = f[400] && f[376] && !f[659] && f[295]; // c2t542i54
	assign leaf[788] = f[400] && f[376] && f[659] && !f[547]; // c2t542i54
	assign leaf[789] = f[400] && f[376] && f[659] && f[547]; // c2t542i54
	assign leaf[790] = !f[378] && !f[400] && !f[425] && !f[149]; // c2t552i55
	assign leaf[791] = !f[378] && !f[400] && !f[425] && f[149]; // c2t552i55
	assign leaf[792] = !f[378] && !f[400] && f[425] && !f[433]; // c2t552i55
	assign leaf[793] = !f[378] && !f[400] && f[425] && f[433]; // c2t552i55
	assign leaf[794] = !f[378] && f[400] && !f[404] && !f[456]; // c2t552i55
	assign leaf[795] = !f[378] && f[400] && !f[404] && f[456]; // c2t552i55
	assign leaf[796] = !f[378] && f[400] && f[404] && !f[343]; // c2t552i55
	assign leaf[797] = !f[378] && f[400] && f[404] && f[343]; // c2t552i55
	assign leaf[798] = f[378] && !f[484] && !f[516] && !f[426]; // c2t552i55
	assign leaf[799] = f[378] && !f[484] && !f[516] && f[426]; // c2t552i55
	assign leaf[800] = f[378] && !f[484] && f[516] && !f[579]; // c2t552i55
	assign leaf[801] = f[378] && !f[484] && f[516] && f[579]; // c2t552i55
	assign leaf[802] = f[378] && f[484] && !f[690] && !f[314]; // c2t552i55
	assign leaf[803] = f[378] && f[484] && !f[690] && f[314]; // c2t552i55
	assign leaf[804] = f[378] && f[484] && f[690]; // c2t552i55
	assign leaf[805] = !f[418] && !f[411] && !f[329] && !f[378]; // c2t562i56
	assign leaf[806] = !f[418] && !f[411] && !f[329] && f[378]; // c2t562i56
	assign leaf[807] = !f[418] && !f[411] && f[329] && !f[324]; // c2t562i56
	assign leaf[808] = !f[418] && !f[411] && f[329] && f[324]; // c2t562i56
	assign leaf[809] = !f[418] && f[411] && !f[353] && !f[540]; // c2t562i56
	assign leaf[810] = !f[418] && f[411] && !f[353] && f[540]; // c2t562i56
	assign leaf[811] = !f[418] && f[411] && f[353] && !f[519]; // c2t562i56
	assign leaf[812] = !f[418] && f[411] && f[353] && f[519]; // c2t562i56
	assign leaf[813] = f[418]; // c2t562i56
	assign leaf[814] = !f[513] && !f[404] && !f[568] && !f[458]; // c2t572i57
	assign leaf[815] = !f[513] && !f[404] && !f[568] && f[458]; // c2t572i57
	assign leaf[816] = !f[513] && !f[404] && f[568] && !f[320]; // c2t572i57
	assign leaf[817] = !f[513] && !f[404] && f[568] && f[320]; // c2t572i57
	assign leaf[818] = !f[513] && f[404] && !f[455] && !f[97]; // c2t572i57
	assign leaf[819] = !f[513] && f[404] && !f[455] && f[97]; // c2t572i57
	assign leaf[820] = !f[513] && f[404] && f[455] && !f[401]; // c2t572i57
	assign leaf[821] = !f[513] && f[404] && f[455] && f[401]; // c2t572i57
	assign leaf[822] = f[513] && !f[459] && !f[351] && !f[552]; // c2t572i57
	assign leaf[823] = f[513] && !f[459] && !f[351] && f[552]; // c2t572i57
	assign leaf[824] = f[513] && !f[459] && f[351] && !f[430]; // c2t572i57
	assign leaf[825] = f[513] && !f[459] && f[351] && f[430]; // c2t572i57
	assign leaf[826] = f[513] && f[459] && !f[294] && !f[186]; // c2t572i57
	assign leaf[827] = f[513] && f[459] && !f[294] && f[186]; // c2t572i57
	assign leaf[828] = f[513] && f[459] && f[294] && !f[96]; // c2t572i57
	assign leaf[829] = f[513] && f[459] && f[294] && f[96]; // c2t572i57
	assign leaf[830] = !f[104] && !f[545] && !f[660] && !f[469]; // c2t582i58
	assign leaf[831] = !f[104] && !f[545] && !f[660] && f[469]; // c2t582i58
	assign leaf[832] = !f[104] && !f[545] && f[660] && !f[464]; // c2t582i58
	assign leaf[833] = !f[104] && !f[545] && f[660] && f[464]; // c2t582i58
	assign leaf[834] = !f[104] && f[545] && !f[427] && !f[343]; // c2t582i58
	assign leaf[835] = !f[104] && f[545] && !f[427] && f[343]; // c2t582i58
	assign leaf[836] = !f[104] && f[545] && f[427] && !f[289]; // c2t582i58
	assign leaf[837] = !f[104] && f[545] && f[427] && f[289]; // c2t582i58
	assign leaf[838] = f[104] && !f[432] && !f[324]; // c2t582i58
	assign leaf[839] = f[104] && !f[432] && f[324]; // c2t582i58
	assign leaf[840] = f[104] && f[432] && !f[593]; // c2t582i58
	assign leaf[841] = f[104] && f[432] && f[593]; // c2t582i58
	assign leaf[842] = !f[677] && !f[622] && !f[219] && !f[103]; // c2t592i59
	assign leaf[843] = !f[677] && !f[622] && !f[219] && f[103]; // c2t592i59
	assign leaf[844] = !f[677] && !f[622] && f[219] && !f[374]; // c2t592i59
	assign leaf[845] = !f[677] && !f[622] && f[219] && f[374]; // c2t592i59
	assign leaf[846] = !f[677] && f[622] && !f[236] && !f[495]; // c2t592i59
	assign leaf[847] = !f[677] && f[622] && !f[236] && f[495]; // c2t592i59
	assign leaf[848] = !f[677] && f[622] && f[236] && !f[661]; // c2t592i59
	assign leaf[849] = !f[677] && f[622] && f[236] && f[661]; // c2t592i59
	assign leaf[850] = f[677] && !f[188]; // c2t592i59
	assign leaf[851] = f[677] && f[188]; // c2t592i59
	assign leaf[852] = !f[513] && !f[404] && !f[257] && !f[571]; // c2t602i60
	assign leaf[853] = !f[513] && !f[404] && !f[257] && f[571]; // c2t602i60
	assign leaf[854] = !f[513] && !f[404] && f[257] && !f[204]; // c2t602i60
	assign leaf[855] = !f[513] && !f[404] && f[257] && f[204]; // c2t602i60
	assign leaf[856] = !f[513] && f[404] && !f[483] && !f[241]; // c2t602i60
	assign leaf[857] = !f[513] && f[404] && !f[483] && f[241]; // c2t602i60
	assign leaf[858] = !f[513] && f[404] && f[483] && !f[401]; // c2t602i60
	assign leaf[859] = !f[513] && f[404] && f[483] && f[401]; // c2t602i60
	assign leaf[860] = f[513] && !f[433] && !f[381] && !f[454]; // c2t602i60
	assign leaf[861] = f[513] && !f[433] && !f[381] && f[454]; // c2t602i60
	assign leaf[862] = f[513] && !f[433] && f[381] && !f[295]; // c2t602i60
	assign leaf[863] = f[513] && !f[433] && f[381] && f[295]; // c2t602i60
	assign leaf[864] = f[513] && f[433] && !f[257] && !f[322]; // c2t602i60
	assign leaf[865] = f[513] && f[433] && !f[257] && f[322]; // c2t602i60
	assign leaf[866] = f[513] && f[433] && f[257] && !f[262]; // c2t602i60
	assign leaf[867] = f[513] && f[433] && f[257] && f[262]; // c2t602i60
	assign leaf[868] = !f[351] && !f[547] && !f[261] && !f[681]; // c2t612i61
	assign leaf[869] = !f[351] && !f[547] && !f[261] && f[681]; // c2t612i61
	assign leaf[870] = !f[351] && !f[547] && f[261] && !f[657]; // c2t612i61
	assign leaf[871] = !f[351] && !f[547] && f[261] && f[657]; // c2t612i61
	assign leaf[872] = !f[351] && f[547] && !f[407] && !f[512]; // c2t612i61
	assign leaf[873] = !f[351] && f[547] && !f[407] && f[512]; // c2t612i61
	assign leaf[874] = !f[351] && f[547] && f[407] && !f[630]; // c2t612i61
	assign leaf[875] = !f[351] && f[547] && f[407] && f[630]; // c2t612i61
	assign leaf[876] = f[351] && !f[437] && !f[605] && !f[524]; // c2t612i61
	assign leaf[877] = f[351] && !f[437] && !f[605] && f[524]; // c2t612i61
	assign leaf[878] = f[351] && !f[437] && f[605] && !f[520]; // c2t612i61
	assign leaf[879] = f[351] && !f[437] && f[605] && f[520]; // c2t612i61
	assign leaf[880] = f[351] && f[437] && !f[659] && !f[482]; // c2t612i61
	assign leaf[881] = f[351] && f[437] && !f[659] && f[482]; // c2t612i61
	assign leaf[882] = f[351] && f[437] && f[659] && !f[257]; // c2t612i61
	assign leaf[883] = f[351] && f[437] && f[659] && f[257]; // c2t612i61
	assign leaf[884] = !f[121] && !f[497] && !f[607] && !f[689]; // c2t622i62
	assign leaf[885] = !f[121] && !f[497] && !f[607] && f[689]; // c2t622i62
	assign leaf[886] = !f[121] && !f[497] && f[607] && !f[551]; // c2t622i62
	assign leaf[887] = !f[121] && !f[497] && f[607] && f[551]; // c2t622i62
	assign leaf[888] = !f[121] && f[497] && !f[633] && !f[609]; // c2t622i62
	assign leaf[889] = !f[121] && f[497] && !f[633] && f[609]; // c2t622i62
	assign leaf[890] = !f[121] && f[497] && f[633] && !f[353]; // c2t622i62
	assign leaf[891] = !f[121] && f[497] && f[633] && f[353]; // c2t622i62
	assign leaf[892] = f[121] && !f[232] && !f[605]; // c2t622i62
	assign leaf[893] = f[121] && !f[232] && f[605] && !f[608]; // c2t622i62
	assign leaf[894] = f[121] && !f[232] && f[605] && f[608]; // c2t622i62
	assign leaf[895] = f[121] && f[232] && !f[467]; // c2t622i62
	assign leaf[896] = f[121] && f[232] && f[467]; // c2t622i62
	assign leaf[897] = !f[709] && !f[409] && !f[460] && !f[494]; // c2t632i63
	assign leaf[898] = !f[709] && !f[409] && !f[460] && f[494]; // c2t632i63
	assign leaf[899] = !f[709] && !f[409] && f[460] && !f[374]; // c2t632i63
	assign leaf[900] = !f[709] && !f[409] && f[460] && f[374]; // c2t632i63
	assign leaf[901] = !f[709] && f[409] && !f[463] && !f[491]; // c2t632i63
	assign leaf[902] = !f[709] && f[409] && !f[463] && f[491]; // c2t632i63
	assign leaf[903] = !f[709] && f[409] && f[463] && !f[679]; // c2t632i63
	assign leaf[904] = !f[709] && f[409] && f[463] && f[679]; // c2t632i63
	assign leaf[905] = f[709]; // c2t632i63
	assign leaf[906] = !f[515] && !f[378] && !f[373] && !f[342]; // c2t642i64
	assign leaf[907] = !f[515] && !f[378] && !f[373] && f[342]; // c2t642i64
	assign leaf[908] = !f[515] && !f[378] && f[373] && !f[154]; // c2t642i64
	assign leaf[909] = !f[515] && !f[378] && f[373] && f[154]; // c2t642i64
	assign leaf[910] = !f[515] && f[378] && !f[175] && !f[212]; // c2t642i64
	assign leaf[911] = !f[515] && f[378] && !f[175] && f[212]; // c2t642i64
	assign leaf[912] = !f[515] && f[378] && f[175] && !f[259]; // c2t642i64
	assign leaf[913] = !f[515] && f[378] && f[175] && f[259]; // c2t642i64
	assign leaf[914] = f[515] && !f[466] && !f[578] && !f[661]; // c2t642i64
	assign leaf[915] = f[515] && !f[466] && !f[578] && f[661]; // c2t642i64
	assign leaf[916] = f[515] && !f[466] && f[578] && !f[597]; // c2t642i64
	assign leaf[917] = f[515] && !f[466] && f[578] && f[597]; // c2t642i64
	assign leaf[918] = f[515] && f[466] && !f[632] && !f[290]; // c2t642i64
	assign leaf[919] = f[515] && f[466] && !f[632] && f[290]; // c2t642i64
	assign leaf[920] = f[515] && f[466] && f[632] && !f[329]; // c2t642i64
	assign leaf[921] = f[515] && f[466] && f[632] && f[329]; // c2t642i64
	assign leaf[922] = !f[154] && !f[133] && !f[219] && !f[213]; // c2t652i65
	assign leaf[923] = !f[154] && !f[133] && !f[219] && f[213]; // c2t652i65
	assign leaf[924] = !f[154] && !f[133] && f[219] && !f[603]; // c2t652i65
	assign leaf[925] = !f[154] && !f[133] && f[219] && f[603]; // c2t652i65
	assign leaf[926] = !f[154] && f[133] && !f[156]; // c2t652i65
	assign leaf[927] = !f[154] && f[133] && f[156] && !f[351]; // c2t652i65
	assign leaf[928] = !f[154] && f[133] && f[156] && f[351]; // c2t652i65
	assign leaf[929] = f[154] && !f[625] && !f[290] && !f[486]; // c2t652i65
	assign leaf[930] = f[154] && !f[625] && !f[290] && f[486]; // c2t652i65
	assign leaf[931] = f[154] && !f[625] && f[290] && !f[299]; // c2t652i65
	assign leaf[932] = f[154] && !f[625] && f[290] && f[299]; // c2t652i65
	assign leaf[933] = f[154] && f[625] && !f[594] && !f[270]; // c2t652i65
	assign leaf[934] = f[154] && f[625] && !f[594] && f[270]; // c2t652i65
	assign leaf[935] = f[154] && f[625] && f[594] && !f[346]; // c2t652i65
	assign leaf[936] = f[154] && f[625] && f[594] && f[346]; // c2t652i65
	assign leaf[937] = !f[242] && !f[183] && !f[326] && !f[240]; // c2t662i66
	assign leaf[938] = !f[242] && !f[183] && !f[326] && f[240]; // c2t662i66
	assign leaf[939] = !f[242] && !f[183] && f[326] && !f[269]; // c2t662i66
	assign leaf[940] = !f[242] && !f[183] && f[326] && f[269]; // c2t662i66
	assign leaf[941] = !f[242] && f[183] && !f[240] && !f[188]; // c2t662i66
	assign leaf[942] = !f[242] && f[183] && !f[240] && f[188]; // c2t662i66
	assign leaf[943] = !f[242] && f[183] && f[240] && !f[500]; // c2t662i66
	assign leaf[944] = !f[242] && f[183] && f[240] && f[500]; // c2t662i66
	assign leaf[945] = f[242] && !f[184] && !f[129] && !f[324]; // c2t662i66
	assign leaf[946] = f[242] && !f[184] && !f[129] && f[324]; // c2t662i66
	assign leaf[947] = f[242] && !f[184] && f[129] && !f[238]; // c2t662i66
	assign leaf[948] = f[242] && !f[184] && f[129] && f[238]; // c2t662i66
	assign leaf[949] = f[242] && f[184] && !f[540] && !f[688]; // c2t662i66
	assign leaf[950] = f[242] && f[184] && !f[540] && f[688]; // c2t662i66
	assign leaf[951] = f[242] && f[184] && f[540] && !f[651]; // c2t662i66
	assign leaf[952] = f[242] && f[184] && f[540] && f[651]; // c2t662i66
	assign leaf[953] = !f[485] && !f[403] && !f[512] && !f[257]; // c2t672i67
	assign leaf[954] = !f[485] && !f[403] && !f[512] && f[257]; // c2t672i67
	assign leaf[955] = !f[485] && !f[403] && f[512] && !f[459]; // c2t672i67
	assign leaf[956] = !f[485] && !f[403] && f[512] && f[459]; // c2t672i67
	assign leaf[957] = !f[485] && f[403] && !f[428] && !f[122]; // c2t672i67
	assign leaf[958] = !f[485] && f[403] && !f[428] && f[122]; // c2t672i67
	assign leaf[959] = !f[485] && f[403] && f[428] && !f[294]; // c2t672i67
	assign leaf[960] = !f[485] && f[403] && f[428] && f[294]; // c2t672i67
	assign leaf[961] = f[485] && !f[690] && !f[685] && !f[433]; // c2t672i67
	assign leaf[962] = f[485] && !f[690] && !f[685] && f[433]; // c2t672i67
	assign leaf[963] = f[485] && !f[690] && f[685] && !f[607]; // c2t672i67
	assign leaf[964] = f[485] && !f[690] && f[685] && f[607]; // c2t672i67
	assign leaf[965] = f[485] && f[690] && !f[187]; // c2t672i67
	assign leaf[966] = f[485] && f[690] && f[187]; // c2t672i67
	assign leaf[967] = !f[323] && !f[261] && !f[292] && !f[399]; // c2t682i68
	assign leaf[968] = !f[323] && !f[261] && !f[292] && f[399]; // c2t682i68
	assign leaf[969] = !f[323] && !f[261] && f[292] && !f[322]; // c2t682i68
	assign leaf[970] = !f[323] && !f[261] && f[292] && f[322]; // c2t682i68
	assign leaf[971] = !f[323] && f[261] && !f[285] && !f[625]; // c2t682i68
	assign leaf[972] = !f[323] && f[261] && !f[285] && f[625]; // c2t682i68
	assign leaf[973] = !f[323] && f[261] && f[285] && !f[484]; // c2t682i68
	assign leaf[974] = !f[323] && f[261] && f[285] && f[484]; // c2t682i68
	assign leaf[975] = f[323] && !f[217] && !f[528] && !f[439]; // c2t682i68
	assign leaf[976] = f[323] && !f[217] && !f[528] && f[439]; // c2t682i68
	assign leaf[977] = f[323] && !f[217] && f[528] && !f[567]; // c2t682i68
	assign leaf[978] = f[323] && !f[217] && f[528] && f[567]; // c2t682i68
	assign leaf[979] = f[323] && f[217] && !f[607] && !f[508]; // c2t682i68
	assign leaf[980] = f[323] && f[217] && !f[607] && f[508]; // c2t682i68
	assign leaf[981] = f[323] && f[217] && f[607] && !f[511]; // c2t682i68
	assign leaf[982] = f[323] && f[217] && f[607] && f[511]; // c2t682i68
	assign leaf[983] = !f[570] && !f[480] && !f[525] && !f[415]; // c2t692i69
	assign leaf[984] = !f[570] && !f[480] && !f[525] && f[415]; // c2t692i69
	assign leaf[985] = !f[570] && !f[480] && f[525] && !f[607]; // c2t692i69
	assign leaf[986] = !f[570] && !f[480] && f[525] && f[607]; // c2t692i69
	assign leaf[987] = !f[570] && f[480] && !f[459]; // c2t692i69
	assign leaf[988] = !f[570] && f[480] && f[459] && !f[440]; // c2t692i69
	assign leaf[989] = !f[570] && f[480] && f[459] && f[440]; // c2t692i69
	assign leaf[990] = f[570] && !f[453] && !f[485] && !f[568]; // c2t692i69
	assign leaf[991] = f[570] && !f[453] && !f[485] && f[568]; // c2t692i69
	assign leaf[992] = f[570] && !f[453] && f[485] && !f[400]; // c2t692i69
	assign leaf[993] = f[570] && !f[453] && f[485] && f[400]; // c2t692i69
	assign leaf[994] = f[570] && f[453] && !f[401] && !f[457]; // c2t692i69
	assign leaf[995] = f[570] && f[453] && !f[401] && f[457]; // c2t692i69
	assign leaf[996] = f[570] && f[453] && f[401] && !f[319]; // c2t692i69
	assign leaf[997] = f[570] && f[453] && f[401] && f[319]; // c2t692i69
	assign leaf[998] = !f[104] && !f[546] && !f[602] && !f[101]; // c2t702i70
	assign leaf[999] = !f[104] && !f[546] && !f[602] && f[101]; // c2t702i70
	assign leaf[1000] = !f[104] && !f[546] && f[602] && !f[492]; // c2t702i70
	assign leaf[1001] = !f[104] && !f[546] && f[602] && f[492]; // c2t702i70
	assign leaf[1002] = !f[104] && f[546] && !f[216] && !f[102]; // c2t702i70
	assign leaf[1003] = !f[104] && f[546] && !f[216] && f[102]; // c2t702i70
	assign leaf[1004] = !f[104] && f[546] && f[216] && !f[352]; // c2t702i70
	assign leaf[1005] = !f[104] && f[546] && f[216] && f[352]; // c2t702i70
	assign leaf[1006] = f[104] && !f[432]; // c2t702i70
	assign leaf[1007] = f[104] && f[432]; // c2t702i70
	assign leaf[1008] = !f[276] && !f[378] && !f[400] && !f[275]; // c2t712i71
	assign leaf[1009] = !f[276] && !f[378] && !f[400] && f[275]; // c2t712i71
	assign leaf[1010] = !f[276] && !f[378] && f[400] && !f[404]; // c2t712i71
	assign leaf[1011] = !f[276] && !f[378] && f[400] && f[404]; // c2t712i71
	assign leaf[1012] = !f[276] && f[378] && !f[214] && !f[658]; // c2t712i71
	assign leaf[1013] = !f[276] && f[378] && !f[214] && f[658]; // c2t712i71
	assign leaf[1014] = !f[276] && f[378] && f[214] && !f[100]; // c2t712i71
	assign leaf[1015] = !f[276] && f[378] && f[214] && f[100]; // c2t712i71
	assign leaf[1016] = f[276]; // c2t712i71
	assign leaf[1017] = !f[712] && !f[677] && !f[322] && !f[657]; // c2t722i72
	assign leaf[1018] = !f[712] && !f[677] && !f[322] && f[657]; // c2t722i72
	assign leaf[1019] = !f[712] && !f[677] && f[322] && !f[325]; // c2t722i72
	assign leaf[1020] = !f[712] && !f[677] && f[322] && f[325]; // c2t722i72
	assign leaf[1021] = !f[712] && f[677]; // c2t722i72
	assign leaf[1022] = f[712] && !f[406]; // c2t722i72
	assign leaf[1023] = f[712] && f[406]; // c2t722i72
	assign leaf[1024] = !f[219] && !f[514] && !f[460] && !f[715]; // c2t732i73
	assign leaf[1025] = !f[219] && !f[514] && !f[460] && f[715]; // c2t732i73
	assign leaf[1026] = !f[219] && !f[514] && f[460] && !f[509]; // c2t732i73
	assign leaf[1027] = !f[219] && !f[514] && f[460] && f[509]; // c2t732i73
	assign leaf[1028] = !f[219] && f[514] && !f[259] && !f[293]; // c2t732i73
	assign leaf[1029] = !f[219] && f[514] && !f[259] && f[293]; // c2t732i73
	assign leaf[1030] = !f[219] && f[514] && f[259] && !f[455]; // c2t732i73
	assign leaf[1031] = !f[219] && f[514] && f[259] && f[455]; // c2t732i73
	assign leaf[1032] = f[219] && !f[622] && !f[599]; // c2t732i73
	assign leaf[1033] = f[219] && !f[622] && f[599]; // c2t732i73
	assign leaf[1034] = f[219] && f[622] && !f[603]; // c2t732i73
	assign leaf[1035] = f[219] && f[622] && f[603]; // c2t732i73
	assign leaf[1036] = !f[411] && !f[173] && !f[356] && !f[463]; // c2t742i74
	assign leaf[1037] = !f[411] && !f[173] && !f[356] && f[463]; // c2t742i74
	assign leaf[1038] = !f[411] && !f[173] && f[356] && !f[463]; // c2t742i74
	assign leaf[1039] = !f[411] && !f[173] && f[356] && f[463]; // c2t742i74
	assign leaf[1040] = !f[411] && f[173] && !f[258] && !f[544]; // c2t742i74
	assign leaf[1041] = !f[411] && f[173] && !f[258] && f[544]; // c2t742i74
	assign leaf[1042] = !f[411] && f[173] && f[258]; // c2t742i74
	assign leaf[1043] = f[411] && !f[493] && !f[512] && !f[600]; // c2t742i74
	assign leaf[1044] = f[411] && !f[493] && !f[512] && f[600]; // c2t742i74
	assign leaf[1045] = f[411] && !f[493] && f[512] && !f[489]; // c2t742i74
	assign leaf[1046] = f[411] && !f[493] && f[512] && f[489]; // c2t742i74
	assign leaf[1047] = f[411] && f[493] && !f[518] && !f[148]; // c2t742i74
	assign leaf[1048] = f[411] && f[493] && !f[518] && f[148]; // c2t742i74
	assign leaf[1049] = f[411] && f[493] && f[518] && !f[555]; // c2t742i74
	assign leaf[1050] = f[411] && f[493] && f[518] && f[555]; // c2t742i74
	assign leaf[1051] = !f[715] && !f[718] && !f[547] && !f[603]; // c2t752i75
	assign leaf[1052] = !f[715] && !f[718] && !f[547] && f[603]; // c2t752i75
	assign leaf[1053] = !f[715] && !f[718] && f[547] && !f[636]; // c2t752i75
	assign leaf[1054] = !f[715] && !f[718] && f[547] && f[636]; // c2t752i75
	assign leaf[1055] = !f[715] && f[718] && !f[492]; // c2t752i75
	assign leaf[1056] = !f[715] && f[718] && f[492]; // c2t752i75
	assign leaf[1057] = f[715] && !f[576] && !f[717]; // c2t752i75
	assign leaf[1058] = f[715] && !f[576] && f[717]; // c2t752i75
	assign leaf[1059] = f[715] && f[576] && !f[295]; // c2t752i75
	assign leaf[1060] = f[715] && f[576] && f[295]; // c2t752i75
	assign leaf[1061] = !f[258] && !f[636] && !f[553] && !f[470]; // c2t762i76
	assign leaf[1062] = !f[258] && !f[636] && !f[553] && f[470]; // c2t762i76
	assign leaf[1063] = !f[258] && !f[636] && f[553] && !f[607]; // c2t762i76
	assign leaf[1064] = !f[258] && !f[636] && f[553] && f[607]; // c2t762i76
	assign leaf[1065] = !f[258] && f[636] && !f[524] && !f[260]; // c2t762i76
	assign leaf[1066] = !f[258] && f[636] && !f[524] && f[260]; // c2t762i76
	assign leaf[1067] = !f[258] && f[636] && f[524] && !f[577]; // c2t762i76
	assign leaf[1068] = !f[258] && f[636] && f[524] && f[577]; // c2t762i76
	assign leaf[1069] = f[258] && !f[455] && !f[635] && !f[244]; // c2t762i76
	assign leaf[1070] = f[258] && !f[455] && !f[635] && f[244]; // c2t762i76
	assign leaf[1071] = f[258] && !f[455] && f[635] && !f[604]; // c2t762i76
	assign leaf[1072] = f[258] && !f[455] && f[635] && f[604]; // c2t762i76
	assign leaf[1073] = f[258] && f[455]; // c2t762i76
	assign leaf[1074] = !f[125] && !f[546] && !f[657] && !f[688]; // c2t772i77
	assign leaf[1075] = !f[125] && !f[546] && !f[657] && f[688]; // c2t772i77
	assign leaf[1076] = !f[125] && !f[546] && f[657] && !f[376]; // c2t772i77
	assign leaf[1077] = !f[125] && !f[546] && f[657] && f[376]; // c2t772i77
	assign leaf[1078] = !f[125] && f[546] && !f[219] && !f[711]; // c2t772i77
	assign leaf[1079] = !f[125] && f[546] && !f[219] && f[711]; // c2t772i77
	assign leaf[1080] = !f[125] && f[546] && f[219] && !f[564]; // c2t772i77
	assign leaf[1081] = !f[125] && f[546] && f[219] && f[564]; // c2t772i77
	assign leaf[1082] = f[125] && !f[240] && !f[381] && !f[300]; // c2t772i77
	assign leaf[1083] = f[125] && !f[240] && !f[381] && f[300]; // c2t772i77
	assign leaf[1084] = f[125] && !f[240] && f[381] && !f[243]; // c2t772i77
	assign leaf[1085] = f[125] && !f[240] && f[381] && f[243]; // c2t772i77
	assign leaf[1086] = f[125] && f[240] && !f[438] && !f[499]; // c2t772i77
	assign leaf[1087] = f[125] && f[240] && !f[438] && f[499]; // c2t772i77
	assign leaf[1088] = f[125] && f[240] && f[438] && !f[266]; // c2t772i77
	assign leaf[1089] = f[125] && f[240] && f[438] && f[266]; // c2t772i77
	assign leaf[1090] = !f[501] && !f[570] && !f[539] && !f[356]; // c2t782i78
	assign leaf[1091] = !f[501] && !f[570] && !f[539] && f[356]; // c2t782i78
	assign leaf[1092] = !f[501] && !f[570] && f[539] && !f[459]; // c2t782i78
	assign leaf[1093] = !f[501] && !f[570] && f[539] && f[459]; // c2t782i78
	assign leaf[1094] = !f[501] && f[570] && !f[406] && !f[524]; // c2t782i78
	assign leaf[1095] = !f[501] && f[570] && !f[406] && f[524]; // c2t782i78
	assign leaf[1096] = !f[501] && f[570] && f[406] && !f[273]; // c2t782i78
	assign leaf[1097] = !f[501] && f[570] && f[406] && f[273]; // c2t782i78
	assign leaf[1098] = f[501] && !f[322]; // c2t782i78
	assign leaf[1099] = f[501] && f[322]; // c2t782i78
	assign leaf[1100] = !f[622] && !f[216] && !f[102] && !f[633]; // c2t792i79
	assign leaf[1101] = !f[622] && !f[216] && !f[102] && f[633]; // c2t792i79
	assign leaf[1102] = !f[622] && !f[216] && f[102] && !f[601]; // c2t792i79
	assign leaf[1103] = !f[622] && !f[216] && f[102] && f[601]; // c2t792i79
	assign leaf[1104] = !f[622] && f[216] && !f[600] && !f[536]; // c2t792i79
	assign leaf[1105] = !f[622] && f[216] && !f[600] && f[536]; // c2t792i79
	assign leaf[1106] = !f[622] && f[216] && f[600] && !f[662]; // c2t792i79
	assign leaf[1107] = !f[622] && f[216] && f[600] && f[662]; // c2t792i79
	assign leaf[1108] = f[622] && !f[634] && !f[551] && !f[352]; // c2t792i79
	assign leaf[1109] = f[622] && !f[634] && !f[551] && f[352]; // c2t792i79
	assign leaf[1110] = f[622] && !f[634] && f[551] && !f[544]; // c2t792i79
	assign leaf[1111] = f[622] && !f[634] && f[551] && f[544]; // c2t792i79
	assign leaf[1112] = f[622] && f[634] && !f[271]; // c2t792i79
	assign leaf[1113] = f[622] && f[634] && f[271]; // c2t792i79
	assign leaf[1114] = !f[677] && !f[659] && !f[689] && !f[684]; // c2t802i80
	assign leaf[1115] = !f[677] && !f[659] && !f[689] && f[684]; // c2t802i80
	assign leaf[1116] = !f[677] && !f[659] && f[689] && !f[572]; // c2t802i80
	assign leaf[1117] = !f[677] && !f[659] && f[689] && f[572]; // c2t802i80
	assign leaf[1118] = !f[677] && f[659] && !f[465] && !f[269]; // c2t802i80
	assign leaf[1119] = !f[677] && f[659] && !f[465] && f[269]; // c2t802i80
	assign leaf[1120] = !f[677] && f[659] && f[465] && !f[229]; // c2t802i80
	assign leaf[1121] = !f[677] && f[659] && f[465] && f[229]; // c2t802i80
	assign leaf[1122] = f[677]; // c2t802i80
	assign leaf[1123] = !f[486] && !f[433] && !f[545] && !f[494]; // c2t812i81
	assign leaf[1124] = !f[486] && !f[433] && !f[545] && f[494]; // c2t812i81
	assign leaf[1125] = !f[486] && !f[433] && f[545] && !f[652]; // c2t812i81
	assign leaf[1126] = !f[486] && !f[433] && f[545] && f[652]; // c2t812i81
	assign leaf[1127] = !f[486] && f[433] && !f[456] && !f[491]; // c2t812i81
	assign leaf[1128] = !f[486] && f[433] && !f[456] && f[491]; // c2t812i81
	assign leaf[1129] = !f[486] && f[433] && f[456] && !f[325]; // c2t812i81
	assign leaf[1130] = !f[486] && f[433] && f[456] && f[325]; // c2t812i81
	assign leaf[1131] = f[486] && !f[432] && !f[324] && !f[568]; // c2t812i81
	assign leaf[1132] = f[486] && !f[432] && !f[324] && f[568]; // c2t812i81
	assign leaf[1133] = f[486] && !f[432] && f[324] && !f[601]; // c2t812i81
	assign leaf[1134] = f[486] && !f[432] && f[324] && f[601]; // c2t812i81
	assign leaf[1135] = f[486] && f[432] && !f[207] && !f[322]; // c2t812i81
	assign leaf[1136] = f[486] && f[432] && !f[207] && f[322]; // c2t812i81
	assign leaf[1137] = f[486] && f[432] && f[207] && !f[567]; // c2t812i81
	assign leaf[1138] = f[486] && f[432] && f[207] && f[567]; // c2t812i81
	assign leaf[1139] = !f[121] && !f[528] && !f[500] && !f[388]; // c2t822i82
	assign leaf[1140] = !f[121] && !f[528] && !f[500] && f[388]; // c2t822i82
	assign leaf[1141] = !f[121] && !f[528] && f[500] && !f[241]; // c2t822i82
	assign leaf[1142] = !f[121] && !f[528] && f[500] && f[241]; // c2t822i82
	assign leaf[1143] = !f[121] && f[528] && !f[500] && !f[512]; // c2t822i82
	assign leaf[1144] = !f[121] && f[528] && !f[500] && f[512]; // c2t822i82
	assign leaf[1145] = !f[121] && f[528] && f[500] && !f[319]; // c2t822i82
	assign leaf[1146] = !f[121] && f[528] && f[500] && f[319]; // c2t822i82
	assign leaf[1147] = f[121] && !f[289] && !f[633] && !f[605]; // c2t822i82
	assign leaf[1148] = f[121] && !f[289] && !f[633] && f[605]; // c2t822i82
	assign leaf[1149] = f[121] && !f[289] && f[633] && !f[498]; // c2t822i82
	assign leaf[1150] = f[121] && !f[289] && f[633] && f[498]; // c2t822i82
	assign leaf[1151] = f[121] && f[289]; // c2t822i82
	assign leaf[1152] = !f[154] && !f[99] && !f[377] && !f[372]; // c2t832i83
	assign leaf[1153] = !f[154] && !f[99] && !f[377] && f[372]; // c2t832i83
	assign leaf[1154] = !f[154] && !f[99] && f[377] && !f[484]; // c2t832i83
	assign leaf[1155] = !f[154] && !f[99] && f[377] && f[484]; // c2t832i83
	assign leaf[1156] = !f[154] && f[99] && !f[566] && !f[487]; // c2t832i83
	assign leaf[1157] = !f[154] && f[99] && !f[566] && f[487]; // c2t832i83
	assign leaf[1158] = !f[154] && f[99] && f[566]; // c2t832i83
	assign leaf[1159] = f[154] && !f[636] && !f[294] && !f[625]; // c2t832i83
	assign leaf[1160] = f[154] && !f[636] && !f[294] && f[625]; // c2t832i83
	assign leaf[1161] = f[154] && !f[636] && f[294] && !f[553]; // c2t832i83
	assign leaf[1162] = f[154] && !f[636] && f[294] && f[553]; // c2t832i83
	assign leaf[1163] = f[154] && f[636] && !f[524] && !f[526]; // c2t832i83
	assign leaf[1164] = f[154] && f[636] && !f[524] && f[526]; // c2t832i83
	assign leaf[1165] = f[154] && f[636] && f[524] && !f[662]; // c2t832i83
	assign leaf[1166] = f[154] && f[636] && f[524] && f[662]; // c2t832i83
	assign leaf[1167] = !f[417] && !f[351] && !f[355] && !f[228]; // c2t842i84
	assign leaf[1168] = !f[417] && !f[351] && !f[355] && f[228]; // c2t842i84
	assign leaf[1169] = !f[417] && !f[351] && f[355] && !f[384]; // c2t842i84
	assign leaf[1170] = !f[417] && !f[351] && f[355] && f[384]; // c2t842i84
	assign leaf[1171] = !f[417] && f[351] && !f[606] && !f[216]; // c2t842i84
	assign leaf[1172] = !f[417] && f[351] && !f[606] && f[216]; // c2t842i84
	assign leaf[1173] = !f[417] && f[351] && f[606] && !f[205]; // c2t842i84
	assign leaf[1174] = !f[417] && f[351] && f[606] && f[205]; // c2t842i84
	assign leaf[1175] = f[417] && !f[240]; // c2t842i84
	assign leaf[1176] = f[417] && f[240]; // c2t842i84
	assign leaf[1177] = !f[709] && !f[712] && !f[134] && !f[104]; // c2t852i85
	assign leaf[1178] = !f[709] && !f[712] && !f[134] && f[104]; // c2t852i85
	assign leaf[1179] = !f[709] && !f[712] && f[134] && !f[273]; // c2t852i85
	assign leaf[1180] = !f[709] && !f[712] && f[134] && f[273]; // c2t852i85
	assign leaf[1181] = !f[709] && f[712]; // c2t852i85
	assign leaf[1182] = f[709]; // c2t852i85
	assign leaf[1183] = !f[374] && !f[125] && !f[209] && !f[326]; // c2t862i86
	assign leaf[1184] = !f[374] && !f[125] && !f[209] && f[326]; // c2t862i86
	assign leaf[1185] = !f[374] && !f[125] && f[209] && !f[599]; // c2t862i86
	assign leaf[1186] = !f[374] && !f[125] && f[209] && f[599]; // c2t862i86
	assign leaf[1187] = !f[374] && f[125] && !f[594] && !f[213]; // c2t862i86
	assign leaf[1188] = !f[374] && f[125] && !f[594] && f[213]; // c2t862i86
	assign leaf[1189] = !f[374] && f[125] && f[594] && !f[578]; // c2t862i86
	assign leaf[1190] = !f[374] && f[125] && f[594] && f[578]; // c2t862i86
	assign leaf[1191] = f[374] && !f[398] && !f[127] && !f[470]; // c2t862i86
	assign leaf[1192] = f[374] && !f[398] && !f[127] && f[470]; // c2t862i86
	assign leaf[1193] = f[374] && !f[398] && f[127] && !f[129]; // c2t862i86
	assign leaf[1194] = f[374] && !f[398] && f[127] && f[129]; // c2t862i86
	assign leaf[1195] = f[374] && f[398] && !f[323] && !f[573]; // c2t862i86
	assign leaf[1196] = f[374] && f[398] && !f[323] && f[573]; // c2t862i86
	assign leaf[1197] = f[374] && f[398] && f[323]; // c2t862i86
	assign leaf[1198] = !f[413] && !f[572] && !f[322] && !f[233]; // c2t872i87
	assign leaf[1199] = !f[413] && !f[572] && !f[322] && f[233]; // c2t872i87
	assign leaf[1200] = !f[413] && !f[572] && f[322] && !f[525]; // c2t872i87
	assign leaf[1201] = !f[413] && !f[572] && f[322] && f[525]; // c2t872i87
	assign leaf[1202] = !f[413] && f[572] && !f[406] && !f[540]; // c2t872i87
	assign leaf[1203] = !f[413] && f[572] && !f[406] && f[540]; // c2t872i87
	assign leaf[1204] = !f[413] && f[572] && f[406] && !f[681]; // c2t872i87
	assign leaf[1205] = !f[413] && f[572] && f[406] && f[681]; // c2t872i87
	assign leaf[1206] = f[413] && !f[464] && !f[174] && !f[624]; // c2t872i87
	assign leaf[1207] = f[413] && !f[464] && !f[174] && f[624]; // c2t872i87
	assign leaf[1208] = f[413] && !f[464] && f[174]; // c2t872i87
	assign leaf[1209] = f[413] && f[464] && !f[490] && !f[212]; // c2t872i87
	assign leaf[1210] = f[413] && f[464] && !f[490] && f[212]; // c2t872i87
	assign leaf[1211] = f[413] && f[464] && f[490] && !f[242]; // c2t872i87
	assign leaf[1212] = f[413] && f[464] && f[490] && f[242]; // c2t872i87
	assign leaf[1213] = !f[486] && !f[432] && !f[209] && !f[492]; // c2t882i88
	assign leaf[1214] = !f[486] && !f[432] && !f[209] && f[492]; // c2t882i88
	assign leaf[1215] = !f[486] && !f[432] && f[209] && !f[568]; // c2t882i88
	assign leaf[1216] = !f[486] && !f[432] && f[209] && f[568]; // c2t882i88
	assign leaf[1217] = !f[486] && f[432] && !f[456] && !f[436]; // c2t882i88
	assign leaf[1218] = !f[486] && f[432] && !f[456] && f[436]; // c2t882i88
	assign leaf[1219] = !f[486] && f[432] && f[456] && !f[325]; // c2t882i88
	assign leaf[1220] = !f[486] && f[432] && f[456] && f[325]; // c2t882i88
	assign leaf[1221] = f[486] && !f[687] && !f[432] && !f[230]; // c2t882i88
	assign leaf[1222] = f[486] && !f[687] && !f[432] && f[230]; // c2t882i88
	assign leaf[1223] = f[486] && !f[687] && f[432] && !f[465]; // c2t882i88
	assign leaf[1224] = f[486] && !f[687] && f[432] && f[465]; // c2t882i88
	assign leaf[1225] = f[486] && f[687] && !f[548] && !f[690]; // c2t882i88
	assign leaf[1226] = f[486] && f[687] && !f[548] && f[690]; // c2t882i88
	assign leaf[1227] = f[486] && f[687] && f[548]; // c2t882i88
	assign leaf[1228] = !f[679] && !f[369] && !f[425] && !f[401]; // c2t892i89
	assign leaf[1229] = !f[679] && !f[369] && !f[425] && f[401]; // c2t892i89
	assign leaf[1230] = !f[679] && !f[369] && f[425] && !f[401]; // c2t892i89
	assign leaf[1231] = !f[679] && !f[369] && f[425] && f[401]; // c2t892i89
	assign leaf[1232] = !f[679] && f[369] && !f[490]; // c2t892i89
	assign leaf[1233] = !f[679] && f[369] && f[490] && !f[440]; // c2t892i89
	assign leaf[1234] = !f[679] && f[369] && f[490] && f[440]; // c2t892i89
	assign leaf[1235] = f[679] && !f[568] && !f[232]; // c2t892i89
	assign leaf[1236] = f[679] && !f[568] && f[232]; // c2t892i89
	assign leaf[1237] = f[679] && f[568] && !f[189]; // c2t892i89
	assign leaf[1238] = f[679] && f[568] && f[189]; // c2t892i89
	assign leaf[1239] = !f[570] && !f[480] && !f[268] && !f[180]; // c2t902i90
	assign leaf[1240] = !f[570] && !f[480] && !f[268] && f[180]; // c2t902i90
	assign leaf[1241] = !f[570] && !f[480] && f[268] && !f[458]; // c2t902i90
	assign leaf[1242] = !f[570] && !f[480] && f[268] && f[458]; // c2t902i90
	assign leaf[1243] = !f[570] && f[480] && !f[461]; // c2t902i90
	assign leaf[1244] = !f[570] && f[480] && f[461]; // c2t902i90
	assign leaf[1245] = f[570] && !f[655] && !f[489] && !f[458]; // c2t902i90
	assign leaf[1246] = f[570] && !f[655] && !f[489] && f[458]; // c2t902i90
	assign leaf[1247] = f[570] && !f[655] && f[489] && !f[681]; // c2t902i90
	assign leaf[1248] = f[570] && !f[655] && f[489] && f[681]; // c2t902i90
	assign leaf[1249] = f[570] && f[655] && !f[403] && !f[406]; // c2t902i90
	assign leaf[1250] = f[570] && f[655] && !f[403] && f[406]; // c2t902i90
	assign leaf[1251] = f[570] && f[655] && f[403] && !f[484]; // c2t902i90
	assign leaf[1252] = f[570] && f[655] && f[403] && f[484]; // c2t902i90
	assign leaf[1253] = !f[512] && !f[575] && !f[714] && !f[654]; // c2t912i91
	assign leaf[1254] = !f[512] && !f[575] && !f[714] && f[654]; // c2t912i91
	assign leaf[1255] = !f[512] && !f[575] && f[714]; // c2t912i91
	assign leaf[1256] = !f[512] && f[575] && !f[403] && !f[100]; // c2t912i91
	assign leaf[1257] = !f[512] && f[575] && !f[403] && f[100]; // c2t912i91
	assign leaf[1258] = !f[512] && f[575] && f[403] && !f[427]; // c2t912i91
	assign leaf[1259] = !f[512] && f[575] && f[403] && f[427]; // c2t912i91
	assign leaf[1260] = f[512] && !f[433] && !f[233] && !f[265]; // c2t912i91
	assign leaf[1261] = f[512] && !f[433] && !f[233] && f[265]; // c2t912i91
	assign leaf[1262] = f[512] && !f[433] && f[233] && !f[595]; // c2t912i91
	assign leaf[1263] = f[512] && !f[433] && f[233] && f[595]; // c2t912i91
	assign leaf[1264] = f[512] && f[433] && !f[457] && !f[186]; // c2t912i91
	assign leaf[1265] = f[512] && f[433] && !f[457] && f[186]; // c2t912i91
	assign leaf[1266] = f[512] && f[433] && f[457] && !f[245]; // c2t912i91
	assign leaf[1267] = f[512] && f[433] && f[457] && f[245]; // c2t912i91
	assign leaf[1268] = !f[455] && !f[611] && !f[430] && !f[346]; // c2t922i92
	assign leaf[1269] = !f[455] && !f[611] && !f[430] && f[346]; // c2t922i92
	assign leaf[1270] = !f[455] && !f[611] && f[430] && !f[484]; // c2t922i92
	assign leaf[1271] = !f[455] && !f[611] && f[430] && f[484]; // c2t922i92
	assign leaf[1272] = !f[455] && f[611] && !f[210]; // c2t922i92
	assign leaf[1273] = !f[455] && f[611] && f[210]; // c2t922i92
	assign leaf[1274] = f[455] && !f[261] && !f[573] && !f[406]; // c2t922i92
	assign leaf[1275] = f[455] && !f[261] && !f[573] && f[406]; // c2t922i92
	assign leaf[1276] = f[455] && !f[261] && f[573] && !f[154]; // c2t922i92
	assign leaf[1277] = f[455] && !f[261] && f[573] && f[154]; // c2t922i92
	assign leaf[1278] = f[455] && f[261] && !f[566] && !f[402]; // c2t922i92
	assign leaf[1279] = f[455] && f[261] && !f[566] && f[402]; // c2t922i92
	assign leaf[1280] = f[455] && f[261] && f[566] && !f[158]; // c2t922i92
	assign leaf[1281] = f[455] && f[261] && f[566] && f[158]; // c2t922i92
	assign leaf[1282] = !f[598] && !f[655] && !f[208] && !f[635]; // c2t932i93
	assign leaf[1283] = !f[598] && !f[655] && !f[208] && f[635]; // c2t932i93
	assign leaf[1284] = !f[598] && !f[655] && f[208] && !f[238]; // c2t932i93
	assign leaf[1285] = !f[598] && !f[655] && f[208] && f[238]; // c2t932i93
	assign leaf[1286] = !f[598] && f[655] && !f[688] && !f[607]; // c2t932i93
	assign leaf[1287] = !f[598] && f[655] && !f[688] && f[607]; // c2t932i93
	assign leaf[1288] = !f[598] && f[655] && f[688]; // c2t932i93
	assign leaf[1289] = f[598] && !f[179] && !f[272] && !f[97]; // c2t932i93
	assign leaf[1290] = f[598] && !f[179] && !f[272] && f[97]; // c2t932i93
	assign leaf[1291] = f[598] && !f[179] && f[272] && !f[264]; // c2t932i93
	assign leaf[1292] = f[598] && !f[179] && f[272] && f[264]; // c2t932i93
	assign leaf[1293] = f[598] && f[179] && !f[268] && !f[409]; // c2t932i93
	assign leaf[1294] = f[598] && f[179] && !f[268] && f[409]; // c2t932i93
	assign leaf[1295] = f[598] && f[179] && f[268] && !f[432]; // c2t932i93
	assign leaf[1296] = f[598] && f[179] && f[268] && f[432]; // c2t932i93
	assign leaf[1297] = !f[397] && !f[154] && !f[374] && !f[493]; // c2t942i94
	assign leaf[1298] = !f[397] && !f[154] && !f[374] && f[493]; // c2t942i94
	assign leaf[1299] = !f[397] && !f[154] && f[374] && !f[182]; // c2t942i94
	assign leaf[1300] = !f[397] && !f[154] && f[374] && f[182]; // c2t942i94
	assign leaf[1301] = !f[397] && f[154] && !f[628] && !f[432]; // c2t942i94
	assign leaf[1302] = !f[397] && f[154] && !f[628] && f[432]; // c2t942i94
	assign leaf[1303] = !f[397] && f[154] && f[628] && !f[266]; // c2t942i94
	assign leaf[1304] = !f[397] && f[154] && f[628] && f[266]; // c2t942i94
	assign leaf[1305] = f[397] && !f[426] && !f[435]; // c2t942i94
	assign leaf[1306] = f[397] && !f[426] && f[435]; // c2t942i94
	assign leaf[1307] = f[397] && f[426] && !f[375]; // c2t942i94
	assign leaf[1308] = f[397] && f[426] && f[375]; // c2t942i94
	assign leaf[1309] = !f[513] && !f[259] && !f[580] && !f[662]; // c2t952i95
	assign leaf[1310] = !f[513] && !f[259] && !f[580] && f[662]; // c2t952i95
	assign leaf[1311] = !f[513] && !f[259] && f[580] && !f[497]; // c2t952i95
	assign leaf[1312] = !f[513] && !f[259] && f[580] && f[497]; // c2t952i95
	assign leaf[1313] = !f[513] && f[259] && !f[579] && !f[428]; // c2t952i95
	assign leaf[1314] = !f[513] && f[259] && !f[579] && f[428]; // c2t952i95
	assign leaf[1315] = !f[513] && f[259] && f[579] && !f[293]; // c2t952i95
	assign leaf[1316] = !f[513] && f[259] && f[579] && f[293]; // c2t952i95
	assign leaf[1317] = f[513] && !f[287] && !f[295] && !f[317]; // c2t952i95
	assign leaf[1318] = f[513] && !f[287] && !f[295] && f[317]; // c2t952i95
	assign leaf[1319] = f[513] && !f[287] && f[295] && !f[431]; // c2t952i95
	assign leaf[1320] = f[513] && !f[287] && f[295] && f[431]; // c2t952i95
	assign leaf[1321] = f[513] && f[287] && !f[595] && !f[579]; // c2t952i95
	assign leaf[1322] = f[513] && f[287] && !f[595] && f[579]; // c2t952i95
	assign leaf[1323] = f[513] && f[287] && f[595]; // c2t952i95
	assign leaf[1324] = !f[715] && !f[121] && !f[570] && !f[296]; // c2t962i96
	assign leaf[1325] = !f[715] && !f[121] && !f[570] && f[296]; // c2t962i96
	assign leaf[1326] = !f[715] && !f[121] && f[570] && !f[400]; // c2t962i96
	assign leaf[1327] = !f[715] && !f[121] && f[570] && f[400]; // c2t962i96
	assign leaf[1328] = !f[715] && f[121] && !f[232] && !f[128]; // c2t962i96
	assign leaf[1329] = !f[715] && f[121] && !f[232] && f[128]; // c2t962i96
	assign leaf[1330] = !f[715] && f[121] && f[232]; // c2t962i96
	assign leaf[1331] = f[715] && !f[494] && !f[178]; // c2t962i96
	assign leaf[1332] = f[715] && !f[494] && f[178]; // c2t962i96
	assign leaf[1333] = f[715] && f[494]; // c2t962i96
	assign leaf[1334] = !f[94] && !f[133] && !f[543] && !f[554]; // c2t972i97
	assign leaf[1335] = !f[94] && !f[133] && !f[543] && f[554]; // c2t972i97
	assign leaf[1336] = !f[94] && !f[133] && f[543] && !f[570]; // c2t972i97
	assign leaf[1337] = !f[94] && !f[133] && f[543] && f[570]; // c2t972i97
	assign leaf[1338] = !f[94] && f[133] && !f[273] && !f[574]; // c2t972i97
	assign leaf[1339] = !f[94] && f[133] && !f[273] && f[574]; // c2t972i97
	assign leaf[1340] = !f[94] && f[133] && f[273] && !f[577]; // c2t972i97
	assign leaf[1341] = !f[94] && f[133] && f[273] && f[577]; // c2t972i97
	assign leaf[1342] = f[94] && !f[149]; // c2t972i97
	assign leaf[1343] = f[94] && f[149]; // c2t972i97
	assign leaf[1344] = !f[487] && !f[433] && !f[174] && !f[653]; // c2t982i98
	assign leaf[1345] = !f[487] && !f[433] && !f[174] && f[653]; // c2t982i98
	assign leaf[1346] = !f[487] && !f[433] && f[174] && !f[609]; // c2t982i98
	assign leaf[1347] = !f[487] && !f[433] && f[174] && f[609]; // c2t982i98
	assign leaf[1348] = !f[487] && f[433] && !f[484] && !f[382]; // c2t982i98
	assign leaf[1349] = !f[487] && f[433] && !f[484] && f[382]; // c2t982i98
	assign leaf[1350] = !f[487] && f[433] && f[484] && !f[294]; // c2t982i98
	assign leaf[1351] = !f[487] && f[433] && f[484] && f[294]; // c2t982i98
	assign leaf[1352] = f[487] && !f[630] && !f[547] && !f[653]; // c2t982i98
	assign leaf[1353] = f[487] && !f[630] && !f[547] && f[653]; // c2t982i98
	assign leaf[1354] = f[487] && !f[630] && f[547] && !f[690]; // c2t982i98
	assign leaf[1355] = f[487] && !f[630] && f[547] && f[690]; // c2t982i98
	assign leaf[1356] = f[487] && f[630] && !f[492] && !f[439]; // c2t982i98
	assign leaf[1357] = f[487] && f[630] && !f[492] && f[439]; // c2t982i98
	assign leaf[1358] = f[487] && f[630] && f[492] && !f[385]; // c2t982i98
	assign leaf[1359] = f[487] && f[630] && f[492] && f[385]; // c2t982i98
	assign leaf[1360] = !f[266] && !f[317] && !f[715] && !f[513]; // c2t992i99
	assign leaf[1361] = !f[266] && !f[317] && !f[715] && f[513]; // c2t992i99
	assign leaf[1362] = !f[266] && !f[317] && f[715]; // c2t992i99
	assign leaf[1363] = !f[266] && f[317] && !f[436] && !f[566]; // c2t992i99
	assign leaf[1364] = !f[266] && f[317] && !f[436] && f[566]; // c2t992i99
	assign leaf[1365] = !f[266] && f[317] && f[436] && !f[380]; // c2t992i99
	assign leaf[1366] = !f[266] && f[317] && f[436] && f[380]; // c2t992i99
	assign leaf[1367] = f[266] && !f[542] && !f[408] && !f[488]; // c2t992i99
	assign leaf[1368] = f[266] && !f[542] && !f[408] && f[488]; // c2t992i99
	assign leaf[1369] = f[266] && !f[542] && f[408] && !f[482]; // c2t992i99
	assign leaf[1370] = f[266] && !f[542] && f[408] && f[482]; // c2t992i99
	assign leaf[1371] = f[266] && f[542] && !f[622] && !f[354]; // c2t992i99
	assign leaf[1372] = f[266] && f[542] && !f[622] && f[354]; // c2t992i99
	assign leaf[1373] = f[266] && f[542] && f[622] && !f[518]; // c2t992i99
	assign leaf[1374] = f[266] && f[542] && f[622] && f[518]; // c2t992i99
endmodule

module decision_tree_leaves_3(input logic [0:783] f, output logic [0:1472] leaf);
	assign leaf[0] = !f[350] && !f[378] && !f[322] && !f[428]; // c3t3i0
	assign leaf[1] = !f[350] && !f[378] && !f[322] && f[428]; // c3t3i0
	assign leaf[2] = !f[350] && !f[378] && f[322] && !f[151]; // c3t3i0
	assign leaf[3] = !f[350] && !f[378] && f[322] && f[151]; // c3t3i0
	assign leaf[4] = !f[350] && f[378] && !f[176] && !f[592]; // c3t3i0
	assign leaf[5] = !f[350] && f[378] && !f[176] && f[592]; // c3t3i0
	assign leaf[6] = !f[350] && f[378] && f[176] && !f[543]; // c3t3i0
	assign leaf[7] = !f[350] && f[378] && f[176] && f[543]; // c3t3i0
	assign leaf[8] = f[350] && !f[489] && !f[290] && !f[179]; // c3t3i0
	assign leaf[9] = f[350] && !f[489] && !f[290] && f[179]; // c3t3i0
	assign leaf[10] = f[350] && !f[489] && f[290] && !f[318]; // c3t3i0
	assign leaf[11] = f[350] && !f[489] && f[290] && f[318]; // c3t3i0
	assign leaf[12] = f[350] && f[489] && !f[517] && !f[515]; // c3t3i0
	assign leaf[13] = f[350] && f[489] && !f[517] && f[515]; // c3t3i0
	assign leaf[14] = f[350] && f[489] && f[517] && !f[536]; // c3t3i0
	assign leaf[15] = f[350] && f[489] && f[517] && f[536]; // c3t3i0
	assign leaf[16] = !f[151] && !f[622] && !f[179] && !f[564]; // c3t13i1
	assign leaf[17] = !f[151] && !f[622] && !f[179] && f[564]; // c3t13i1
	assign leaf[18] = !f[151] && !f[622] && f[179] && !f[317]; // c3t13i1
	assign leaf[19] = !f[151] && !f[622] && f[179] && f[317]; // c3t13i1
	assign leaf[20] = !f[151] && f[622] && !f[351] && !f[379]; // c3t13i1
	assign leaf[21] = !f[151] && f[622] && !f[351] && f[379]; // c3t13i1
	assign leaf[22] = !f[151] && f[622] && f[351] && !f[486]; // c3t13i1
	assign leaf[23] = !f[151] && f[622] && f[351] && f[486]; // c3t13i1
	assign leaf[24] = f[151] && !f[514] && !f[289] && !f[518]; // c3t13i1
	assign leaf[25] = f[151] && !f[514] && !f[289] && f[518]; // c3t13i1
	assign leaf[26] = f[151] && !f[514] && f[289] && !f[267]; // c3t13i1
	assign leaf[27] = f[151] && !f[514] && f[289] && f[267]; // c3t13i1
	assign leaf[28] = f[151] && f[514] && !f[321] && !f[679]; // c3t13i1
	assign leaf[29] = f[151] && f[514] && !f[321] && f[679]; // c3t13i1
	assign leaf[30] = f[151] && f[514] && f[321] && !f[459]; // c3t13i1
	assign leaf[31] = f[151] && f[514] && f[321] && f[459]; // c3t13i1
	assign leaf[32] = !f[350] && !f[378] && !f[322] && !f[406]; // c3t23i2
	assign leaf[33] = !f[350] && !f[378] && !f[322] && f[406]; // c3t23i2
	assign leaf[34] = !f[350] && !f[378] && f[322] && !f[153]; // c3t23i2
	assign leaf[35] = !f[350] && !f[378] && f[322] && f[153]; // c3t23i2
	assign leaf[36] = !f[350] && f[378] && !f[318] && !f[543]; // c3t23i2
	assign leaf[37] = !f[350] && f[378] && !f[318] && f[543]; // c3t23i2
	assign leaf[38] = !f[350] && f[378] && f[318] && !f[148]; // c3t23i2
	assign leaf[39] = !f[350] && f[378] && f[318] && f[148]; // c3t23i2
	assign leaf[40] = f[350] && !f[517] && !f[487] && !f[316]; // c3t23i2
	assign leaf[41] = f[350] && !f[517] && !f[487] && f[316]; // c3t23i2
	assign leaf[42] = f[350] && !f[517] && f[487] && !f[542]; // c3t23i2
	assign leaf[43] = f[350] && !f[517] && f[487] && f[542]; // c3t23i2
	assign leaf[44] = f[350] && f[517] && !f[462] && !f[410]; // c3t23i2
	assign leaf[45] = f[350] && f[517] && !f[462] && f[410]; // c3t23i2
	assign leaf[46] = f[350] && f[517] && f[462] && !f[594]; // c3t23i2
	assign leaf[47] = f[350] && f[517] && f[462] && f[594]; // c3t23i2
	assign leaf[48] = !f[490] && !f[317] && !f[487] && !f[291]; // c3t33i3
	assign leaf[49] = !f[490] && !f[317] && !f[487] && f[291]; // c3t33i3
	assign leaf[50] = !f[490] && !f[317] && f[487] && !f[515]; // c3t33i3
	assign leaf[51] = !f[490] && !f[317] && f[487] && f[515]; // c3t33i3
	assign leaf[52] = !f[490] && f[317] && !f[147] && !f[322]; // c3t33i3
	assign leaf[53] = !f[490] && f[317] && !f[147] && f[322]; // c3t33i3
	assign leaf[54] = !f[490] && f[317] && f[147] && !f[259]; // c3t33i3
	assign leaf[55] = !f[490] && f[317] && f[147] && f[259]; // c3t33i3
	assign leaf[56] = f[490] && !f[178] && !f[649] && !f[297]; // c3t33i3
	assign leaf[57] = f[490] && !f[178] && !f[649] && f[297]; // c3t33i3
	assign leaf[58] = f[490] && !f[178] && f[649] && !f[515]; // c3t33i3
	assign leaf[59] = f[490] && !f[178] && f[649] && f[515]; // c3t33i3
	assign leaf[60] = f[490] && f[178] && !f[657] && !f[714]; // c3t33i3
	assign leaf[61] = f[490] && f[178] && !f[657] && f[714]; // c3t33i3
	assign leaf[62] = f[490] && f[178] && f[657] && !f[545]; // c3t33i3
	assign leaf[63] = f[490] && f[178] && f[657] && f[545]; // c3t33i3
	assign leaf[64] = !f[518] && !f[316] && !f[291] && !f[515]; // c3t43i4
	assign leaf[65] = !f[518] && !f[316] && !f[291] && f[515]; // c3t43i4
	assign leaf[66] = !f[518] && !f[316] && f[291] && !f[176]; // c3t43i4
	assign leaf[67] = !f[518] && !f[316] && f[291] && f[176]; // c3t43i4
	assign leaf[68] = !f[518] && f[316] && !f[399] && !f[292]; // c3t43i4
	assign leaf[69] = !f[518] && f[316] && !f[399] && f[292]; // c3t43i4
	assign leaf[70] = !f[518] && f[316] && f[399] && !f[121]; // c3t43i4
	assign leaf[71] = !f[518] && f[316] && f[399] && f[121]; // c3t43i4
	assign leaf[72] = f[518] && !f[624] && !f[463] && !f[352]; // c3t43i4
	assign leaf[73] = f[518] && !f[624] && !f[463] && f[352]; // c3t43i4
	assign leaf[74] = f[518] && !f[624] && f[463] && !f[650]; // c3t43i4
	assign leaf[75] = f[518] && !f[624] && f[463] && f[650]; // c3t43i4
	assign leaf[76] = f[518] && f[624] && !f[351] && !f[203]; // c3t43i4
	assign leaf[77] = f[518] && f[624] && !f[351] && f[203]; // c3t43i4
	assign leaf[78] = f[518] && f[624] && f[351] && !f[485]; // c3t43i4
	assign leaf[79] = f[518] && f[624] && f[351] && f[485]; // c3t43i4
	assign leaf[80] = !f[152] && !f[180] && !f[563] && !f[507]; // c3t53i5
	assign leaf[81] = !f[152] && !f[180] && !f[563] && f[507]; // c3t53i5
	assign leaf[82] = !f[152] && !f[180] && f[563] && !f[482]; // c3t53i5
	assign leaf[83] = !f[152] && !f[180] && f[563] && f[482]; // c3t53i5
	assign leaf[84] = !f[152] && f[180] && !f[317] && !f[515]; // c3t53i5
	assign leaf[85] = !f[152] && f[180] && !f[317] && f[515]; // c3t53i5
	assign leaf[86] = !f[152] && f[180] && f[317] && !f[228]; // c3t53i5
	assign leaf[87] = !f[152] && f[180] && f[317] && f[228]; // c3t53i5
	assign leaf[88] = f[152] && !f[485] && !f[296] && !f[239]; // c3t53i5
	assign leaf[89] = f[152] && !f[485] && !f[296] && f[239]; // c3t53i5
	assign leaf[90] = f[152] && !f[485] && f[296] && !f[516]; // c3t53i5
	assign leaf[91] = f[152] && !f[485] && f[296] && f[516]; // c3t53i5
	assign leaf[92] = f[152] && f[485] && !f[295] && !f[678]; // c3t53i5
	assign leaf[93] = f[152] && f[485] && !f[295] && f[678]; // c3t53i5
	assign leaf[94] = f[152] && f[485] && f[295] && !f[431]; // c3t53i5
	assign leaf[95] = f[152] && f[485] && f[295] && f[431]; // c3t53i5
	assign leaf[96] = !f[490] && !f[343] && !f[485] && !f[263]; // c3t63i6
	assign leaf[97] = !f[490] && !f[343] && !f[485] && f[263]; // c3t63i6
	assign leaf[98] = !f[490] && !f[343] && f[485] && !f[203]; // c3t63i6
	assign leaf[99] = !f[490] && !f[343] && f[485] && f[203]; // c3t63i6
	assign leaf[100] = !f[490] && f[343] && !f[287] && !f[149]; // c3t63i6
	assign leaf[101] = !f[490] && f[343] && !f[287] && f[149]; // c3t63i6
	assign leaf[102] = !f[490] && f[343] && f[287] && !f[289]; // c3t63i6
	assign leaf[103] = !f[490] && f[343] && f[287] && f[289]; // c3t63i6
	assign leaf[104] = f[490] && !f[324] && !f[682] && !f[203]; // c3t63i6
	assign leaf[105] = f[490] && !f[324] && !f[682] && f[203]; // c3t63i6
	assign leaf[106] = f[490] && !f[324] && f[682] && !f[545]; // c3t63i6
	assign leaf[107] = f[490] && !f[324] && f[682] && f[545]; // c3t63i6
	assign leaf[108] = f[490] && f[324] && !f[181] && !f[101]; // c3t63i6
	assign leaf[109] = f[490] && f[324] && !f[181] && f[101]; // c3t63i6
	assign leaf[110] = f[490] && f[324] && f[181] && !f[654]; // c3t63i6
	assign leaf[111] = f[490] && f[324] && f[181] && f[654]; // c3t63i6
	assign leaf[112] = !f[177] && !f[623] && !f[122] && !f[678]; // c3t73i7
	assign leaf[113] = !f[177] && !f[623] && !f[122] && f[678]; // c3t73i7
	assign leaf[114] = !f[177] && !f[623] && f[122] && !f[629]; // c3t73i7
	assign leaf[115] = !f[177] && !f[623] && f[122] && f[629]; // c3t73i7
	assign leaf[116] = !f[177] && f[623] && !f[324] && !f[511]; // c3t73i7
	assign leaf[117] = !f[177] && f[623] && !f[324] && f[511]; // c3t73i7
	assign leaf[118] = !f[177] && f[623] && f[324] && !f[486]; // c3t73i7
	assign leaf[119] = !f[177] && f[623] && f[324] && f[486]; // c3t73i7
	assign leaf[120] = f[177] && !f[288] && !f[657] && !f[320]; // c3t73i7
	assign leaf[121] = f[177] && !f[288] && !f[657] && f[320]; // c3t73i7
	assign leaf[122] = f[177] && !f[288] && f[657] && !f[314]; // c3t73i7
	assign leaf[123] = f[177] && !f[288] && f[657] && f[314]; // c3t73i7
	assign leaf[124] = f[177] && f[288] && !f[264] && !f[344]; // c3t73i7
	assign leaf[125] = f[177] && f[288] && !f[264] && f[344]; // c3t73i7
	assign leaf[126] = f[177] && f[288] && f[264] && !f[371]; // c3t73i7
	assign leaf[127] = f[177] && f[288] && f[264] && f[371]; // c3t73i7
	assign leaf[128] = !f[655] && !f[710] && !f[627] && !f[175]; // c3t83i8
	assign leaf[129] = !f[655] && !f[710] && !f[627] && f[175]; // c3t83i8
	assign leaf[130] = !f[655] && !f[710] && f[627] && !f[457]; // c3t83i8
	assign leaf[131] = !f[655] && !f[710] && f[627] && f[457]; // c3t83i8
	assign leaf[132] = !f[655] && f[710] && !f[485] && !f[265]; // c3t83i8
	assign leaf[133] = !f[655] && f[710] && !f[485] && f[265]; // c3t83i8
	assign leaf[134] = !f[655] && f[710] && f[485]; // c3t83i8
	assign leaf[135] = f[655] && !f[517] && !f[318] && !f[343]; // c3t83i8
	assign leaf[136] = f[655] && !f[517] && !f[318] && f[343]; // c3t83i8
	assign leaf[137] = f[655] && !f[517] && f[318] && !f[148]; // c3t83i8
	assign leaf[138] = f[655] && !f[517] && f[318] && f[148]; // c3t83i8
	assign leaf[139] = f[655] && f[517] && !f[603] && !f[153]; // c3t83i8
	assign leaf[140] = f[655] && f[517] && !f[603] && f[153]; // c3t83i8
	assign leaf[141] = f[655] && f[517] && f[603] && !f[290]; // c3t83i8
	assign leaf[142] = f[655] && f[517] && f[603] && f[290]; // c3t83i8
	assign leaf[143] = !f[518] && !f[344] && !f[516] && !f[485]; // c3t93i9
	assign leaf[144] = !f[518] && !f[344] && !f[516] && f[485]; // c3t93i9
	assign leaf[145] = !f[518] && !f[344] && f[516] && !f[488]; // c3t93i9
	assign leaf[146] = !f[518] && !f[344] && f[516] && f[488]; // c3t93i9
	assign leaf[147] = !f[518] && f[344] && !f[288] && !f[348]; // c3t93i9
	assign leaf[148] = !f[518] && f[344] && !f[288] && f[348]; // c3t93i9
	assign leaf[149] = !f[518] && f[344] && f[288] && !f[291]; // c3t93i9
	assign leaf[150] = !f[518] && f[344] && f[288] && f[291]; // c3t93i9
	assign leaf[151] = f[518] && !f[463] && !f[352] && !f[632]; // c3t93i9
	assign leaf[152] = f[518] && !f[463] && !f[352] && f[632]; // c3t93i9
	assign leaf[153] = f[518] && !f[463] && f[352] && !f[373]; // c3t93i9
	assign leaf[154] = f[518] && !f[463] && f[352] && f[373]; // c3t93i9
	assign leaf[155] = f[518] && f[463] && !f[623] && !f[536]; // c3t93i9
	assign leaf[156] = f[518] && f[463] && !f[623] && f[536]; // c3t93i9
	assign leaf[157] = f[518] && f[463] && f[623] && !f[352]; // c3t93i9
	assign leaf[158] = f[518] && f[463] && f[623] && f[352]; // c3t93i9
	assign leaf[159] = !f[655] && !f[400] && !f[495] && !f[469]; // c3t103i10
	assign leaf[160] = !f[655] && !f[400] && !f[495] && f[469]; // c3t103i10
	assign leaf[161] = !f[655] && !f[400] && f[495] && !f[458]; // c3t103i10
	assign leaf[162] = !f[655] && !f[400] && f[495] && f[458]; // c3t103i10
	assign leaf[163] = !f[655] && f[400] && !f[200] && !f[710]; // c3t103i10
	assign leaf[164] = !f[655] && f[400] && !f[200] && f[710]; // c3t103i10
	assign leaf[165] = !f[655] && f[400] && f[200] && !f[314]; // c3t103i10
	assign leaf[166] = !f[655] && f[400] && f[200] && f[314]; // c3t103i10
	assign leaf[167] = f[655] && !f[291] && !f[544] && !f[317]; // c3t103i10
	assign leaf[168] = f[655] && !f[291] && !f[544] && f[317]; // c3t103i10
	assign leaf[169] = f[655] && !f[291] && f[544] && !f[489]; // c3t103i10
	assign leaf[170] = f[655] && !f[291] && f[544] && f[489]; // c3t103i10
	assign leaf[171] = f[655] && f[291] && !f[149] && !f[319]; // c3t103i10
	assign leaf[172] = f[655] && f[291] && !f[149] && f[319]; // c3t103i10
	assign leaf[173] = f[655] && f[291] && f[149] && !f[261]; // c3t103i10
	assign leaf[174] = f[655] && f[291] && f[149] && f[261]; // c3t103i10
	assign leaf[175] = !f[428] && !f[523] && !f[565] && !f[181]; // c3t113i11
	assign leaf[176] = !f[428] && !f[523] && !f[565] && f[181]; // c3t113i11
	assign leaf[177] = !f[428] && !f[523] && f[565] && !f[353]; // c3t113i11
	assign leaf[178] = !f[428] && !f[523] && f[565] && f[353]; // c3t113i11
	assign leaf[179] = !f[428] && f[523] && !f[240] && !f[243]; // c3t113i11
	assign leaf[180] = !f[428] && f[523] && !f[240] && f[243]; // c3t113i11
	assign leaf[181] = !f[428] && f[523] && f[240] && !f[516]; // c3t113i11
	assign leaf[182] = !f[428] && f[523] && f[240] && f[516]; // c3t113i11
	assign leaf[183] = f[428] && !f[680] && !f[343] && !f[202]; // c3t113i11
	assign leaf[184] = f[428] && !f[680] && !f[343] && f[202]; // c3t113i11
	assign leaf[185] = f[428] && !f[680] && f[343] && !f[318]; // c3t113i11
	assign leaf[186] = f[428] && !f[680] && f[343] && f[318]; // c3t113i11
	assign leaf[187] = f[428] && f[680] && !f[318] && !f[539]; // c3t113i11
	assign leaf[188] = f[428] && f[680] && !f[318] && f[539]; // c3t113i11
	assign leaf[189] = f[428] && f[680] && f[318] && !f[204]; // c3t113i11
	assign leaf[190] = f[428] && f[680] && f[318] && f[204]; // c3t113i11
	assign leaf[191] = !f[371] && !f[291] && !f[182] && !f[578]; // c3t123i12
	assign leaf[192] = !f[371] && !f[291] && !f[182] && f[578]; // c3t123i12
	assign leaf[193] = !f[371] && !f[291] && f[182] && !f[317]; // c3t123i12
	assign leaf[194] = !f[371] && !f[291] && f[182] && f[317]; // c3t123i12
	assign leaf[195] = !f[371] && f[291] && !f[266] && !f[651]; // c3t123i12
	assign leaf[196] = !f[371] && f[291] && !f[266] && f[651]; // c3t123i12
	assign leaf[197] = !f[371] && f[291] && f[266] && !f[123]; // c3t123i12
	assign leaf[198] = !f[371] && f[291] && f[266] && f[123]; // c3t123i12
	assign leaf[199] = f[371] && !f[320] && !f[259] && !f[149]; // c3t123i12
	assign leaf[200] = f[371] && !f[320] && !f[259] && f[149]; // c3t123i12
	assign leaf[201] = f[371] && !f[320] && f[259] && !f[375]; // c3t123i12
	assign leaf[202] = f[371] && !f[320] && f[259] && f[375]; // c3t123i12
	assign leaf[203] = f[371] && f[320] && !f[151] && !f[256]; // c3t123i12
	assign leaf[204] = f[371] && f[320] && !f[151] && f[256]; // c3t123i12
	assign leaf[205] = f[371] && f[320] && f[151] && !f[260]; // c3t123i12
	assign leaf[206] = f[371] && f[320] && f[151] && f[260]; // c3t123i12
	assign leaf[207] = !f[456] && !f[518] && !f[515] && !f[342]; // c3t133i13
	assign leaf[208] = !f[456] && !f[518] && !f[515] && f[342]; // c3t133i13
	assign leaf[209] = !f[456] && !f[518] && f[515] && !f[460]; // c3t133i13
	assign leaf[210] = !f[456] && !f[518] && f[515] && f[460]; // c3t133i13
	assign leaf[211] = !f[456] && f[518] && !f[594] && !f[463]; // c3t133i13
	assign leaf[212] = !f[456] && f[518] && !f[594] && f[463]; // c3t133i13
	assign leaf[213] = !f[456] && f[518] && f[594] && !f[325]; // c3t133i13
	assign leaf[214] = !f[456] && f[518] && f[594] && f[325]; // c3t133i13
	assign leaf[215] = f[456] && !f[678] && !f[351] && !f[633]; // c3t133i13
	assign leaf[216] = f[456] && !f[678] && !f[351] && f[633]; // c3t133i13
	assign leaf[217] = f[456] && !f[678] && f[351] && !f[343]; // c3t133i13
	assign leaf[218] = f[456] && !f[678] && f[351] && f[343]; // c3t133i13
	assign leaf[219] = f[456] && f[678] && !f[292] && !f[322]; // c3t133i13
	assign leaf[220] = f[456] && f[678] && !f[292] && f[322]; // c3t133i13
	assign leaf[221] = f[456] && f[678] && f[292]; // c3t133i13
	assign leaf[222] = !f[351] && !f[546] && !f[294] && !f[682]; // c3t143i14
	assign leaf[223] = !f[351] && !f[546] && !f[294] && f[682]; // c3t143i14
	assign leaf[224] = !f[351] && !f[546] && f[294] && !f[298]; // c3t143i14
	assign leaf[225] = !f[351] && !f[546] && f[294] && f[298]; // c3t143i14
	assign leaf[226] = !f[351] && f[546] && !f[464] && !f[353]; // c3t143i14
	assign leaf[227] = !f[351] && f[546] && !f[464] && f[353]; // c3t143i14
	assign leaf[228] = !f[351] && f[546] && f[464] && !f[678]; // c3t143i14
	assign leaf[229] = !f[351] && f[546] && f[464] && f[678]; // c3t143i14
	assign leaf[230] = f[351] && !f[269] && !f[271] && !f[175]; // c3t143i14
	assign leaf[231] = f[351] && !f[269] && !f[271] && f[175]; // c3t143i14
	assign leaf[232] = f[351] && !f[269] && f[271] && !f[345]; // c3t143i14
	assign leaf[233] = f[351] && !f[269] && f[271] && f[345]; // c3t143i14
	assign leaf[234] = f[351] && f[269] && !f[183] && !f[127]; // c3t143i14
	assign leaf[235] = f[351] && f[269] && !f[183] && f[127]; // c3t143i14
	assign leaf[236] = f[351] && f[269] && f[183] && !f[514]; // c3t143i14
	assign leaf[237] = f[351] && f[269] && f[183] && f[514]; // c3t143i14
	assign leaf[238] = !f[429] && !f[495] && !f[469] && !f[521]; // c3t153i15
	assign leaf[239] = !f[429] && !f[495] && !f[469] && f[521]; // c3t153i15
	assign leaf[240] = !f[429] && !f[495] && f[469] && !f[265]; // c3t153i15
	assign leaf[241] = !f[429] && !f[495] && f[469] && f[265]; // c3t153i15
	assign leaf[242] = !f[429] && f[495] && !f[398] && !f[262]; // c3t153i15
	assign leaf[243] = !f[429] && f[495] && !f[398] && f[262]; // c3t153i15
	assign leaf[244] = !f[429] && f[495] && f[398] && !f[371]; // c3t153i15
	assign leaf[245] = !f[429] && f[495] && f[398] && f[371]; // c3t153i15
	assign leaf[246] = f[429] && !f[511] && !f[318] && !f[343]; // c3t153i15
	assign leaf[247] = f[429] && !f[511] && !f[318] && f[343]; // c3t153i15
	assign leaf[248] = f[429] && !f[511] && f[318] && !f[231]; // c3t153i15
	assign leaf[249] = f[429] && !f[511] && f[318] && f[231]; // c3t153i15
	assign leaf[250] = f[429] && f[511] && !f[453] && !f[456]; // c3t153i15
	assign leaf[251] = f[429] && f[511] && !f[453] && f[456]; // c3t153i15
	assign leaf[252] = f[429] && f[511] && f[453] && !f[464]; // c3t153i15
	assign leaf[253] = f[429] && f[511] && f[453] && f[464]; // c3t153i15
	assign leaf[254] = !f[372] && !f[212] && !f[173] && !f[487]; // c3t163i16
	assign leaf[255] = !f[372] && !f[212] && !f[173] && f[487]; // c3t163i16
	assign leaf[256] = !f[372] && !f[212] && f[173] && !f[493]; // c3t163i16
	assign leaf[257] = !f[372] && !f[212] && f[173] && f[493]; // c3t163i16
	assign leaf[258] = !f[372] && f[212] && !f[319] && !f[405]; // c3t163i16
	assign leaf[259] = !f[372] && f[212] && !f[319] && f[405]; // c3t163i16
	assign leaf[260] = !f[372] && f[212] && f[319] && !f[294]; // c3t163i16
	assign leaf[261] = !f[372] && f[212] && f[319] && f[294]; // c3t163i16
	assign leaf[262] = f[372] && !f[321] && !f[492] && !f[259]; // c3t163i16
	assign leaf[263] = f[372] && !f[321] && !f[492] && f[259]; // c3t163i16
	assign leaf[264] = f[372] && !f[321] && f[492] && !f[650]; // c3t163i16
	assign leaf[265] = f[372] && !f[321] && f[492] && f[650]; // c3t163i16
	assign leaf[266] = f[372] && f[321] && !f[455] && !f[288]; // c3t163i16
	assign leaf[267] = f[372] && f[321] && !f[455] && f[288]; // c3t163i16
	assign leaf[268] = f[372] && f[321] && f[455] && !f[202]; // c3t163i16
	assign leaf[269] = f[372] && f[321] && f[455] && f[202]; // c3t163i16
	assign leaf[270] = !f[427] && !f[202] && !f[292] && !f[317]; // c3t173i17
	assign leaf[271] = !f[427] && !f[202] && !f[292] && f[317]; // c3t173i17
	assign leaf[272] = !f[427] && !f[202] && f[292] && !f[267]; // c3t173i17
	assign leaf[273] = !f[427] && !f[202] && f[292] && f[267]; // c3t173i17
	assign leaf[274] = !f[427] && f[202] && !f[580] && !f[492]; // c3t173i17
	assign leaf[275] = !f[427] && f[202] && !f[580] && f[492]; // c3t173i17
	assign leaf[276] = !f[427] && f[202] && f[580] && !f[237]; // c3t173i17
	assign leaf[277] = !f[427] && f[202] && f[580] && f[237]; // c3t173i17
	assign leaf[278] = f[427] && !f[357] && !f[681] && !f[128]; // c3t173i17
	assign leaf[279] = f[427] && !f[357] && !f[681] && f[128]; // c3t173i17
	assign leaf[280] = f[427] && !f[357] && f[681] && !f[318]; // c3t173i17
	assign leaf[281] = f[427] && !f[357] && f[681] && f[318]; // c3t173i17
	assign leaf[282] = f[427] && f[357] && !f[189] && !f[229]; // c3t173i17
	assign leaf[283] = f[427] && f[357] && !f[189] && f[229]; // c3t173i17
	assign leaf[284] = f[427] && f[357] && f[189] && !f[400]; // c3t173i17
	assign leaf[285] = f[427] && f[357] && f[189] && f[400]; // c3t173i17
	assign leaf[286] = !f[551] && !f[184] && !f[581] && !f[373]; // c3t183i18
	assign leaf[287] = !f[551] && !f[184] && !f[581] && f[373]; // c3t183i18
	assign leaf[288] = !f[551] && !f[184] && f[581] && !f[265]; // c3t183i18
	assign leaf[289] = !f[551] && !f[184] && f[581] && f[265]; // c3t183i18
	assign leaf[290] = !f[551] && f[184] && !f[292] && !f[548]; // c3t183i18
	assign leaf[291] = !f[551] && f[184] && !f[292] && f[548]; // c3t183i18
	assign leaf[292] = !f[551] && f[184] && f[292] && !f[125]; // c3t183i18
	assign leaf[293] = !f[551] && f[184] && f[292] && f[125]; // c3t183i18
	assign leaf[294] = f[551] && !f[371] && !f[239] && !f[291]; // c3t183i18
	assign leaf[295] = f[551] && !f[371] && !f[239] && f[291]; // c3t183i18
	assign leaf[296] = f[551] && !f[371] && f[239] && !f[545]; // c3t183i18
	assign leaf[297] = f[551] && !f[371] && f[239] && f[545]; // c3t183i18
	assign leaf[298] = f[551] && f[371] && !f[347] && !f[400]; // c3t183i18
	assign leaf[299] = f[551] && f[371] && !f[347] && f[400]; // c3t183i18
	assign leaf[300] = f[551] && f[371] && f[347] && !f[482]; // c3t183i18
	assign leaf[301] = f[551] && f[371] && f[347] && f[482]; // c3t183i18
	assign leaf[302] = !f[373] && !f[536] && !f[682] && !f[123]; // c3t193i19
	assign leaf[303] = !f[373] && !f[536] && !f[682] && f[123]; // c3t193i19
	assign leaf[304] = !f[373] && !f[536] && f[682] && !f[570]; // c3t193i19
	assign leaf[305] = !f[373] && !f[536] && f[682] && f[570]; // c3t193i19
	assign leaf[306] = !f[373] && f[536] && !f[327] && !f[429]; // c3t193i19
	assign leaf[307] = !f[373] && f[536] && !f[327] && f[429]; // c3t193i19
	assign leaf[308] = !f[373] && f[536] && f[327] && !f[458]; // c3t193i19
	assign leaf[309] = !f[373] && f[536] && f[327] && f[458]; // c3t193i19
	assign leaf[310] = f[373] && !f[321] && !f[345] && !f[371]; // c3t193i19
	assign leaf[311] = f[373] && !f[321] && !f[345] && f[371]; // c3t193i19
	assign leaf[312] = f[373] && !f[321] && f[345] && !f[200]; // c3t193i19
	assign leaf[313] = f[373] && !f[321] && f[345] && f[200]; // c3t193i19
	assign leaf[314] = f[373] && f[321] && !f[152] && !f[206]; // c3t193i19
	assign leaf[315] = f[373] && f[321] && !f[152] && f[206]; // c3t193i19
	assign leaf[316] = f[373] && f[321] && f[152] && !f[289]; // c3t193i19
	assign leaf[317] = f[373] && f[321] && f[152] && f[289]; // c3t193i19
	assign leaf[318] = !f[578] && !f[457] && !f[625] && !f[679]; // c3t203i20
	assign leaf[319] = !f[578] && !f[457] && !f[625] && f[679]; // c3t203i20
	assign leaf[320] = !f[578] && !f[457] && f[625] && !f[487]; // c3t203i20
	assign leaf[321] = !f[578] && !f[457] && f[625] && f[487]; // c3t203i20
	assign leaf[322] = !f[578] && f[457] && !f[678] && !f[708]; // c3t203i20
	assign leaf[323] = !f[578] && f[457] && !f[678] && f[708]; // c3t203i20
	assign leaf[324] = !f[578] && f[457] && f[678] && !f[511]; // c3t203i20
	assign leaf[325] = !f[578] && f[457] && f[678] && f[511]; // c3t203i20
	assign leaf[326] = f[578] && !f[712] && !f[176] && !f[651]; // c3t203i20
	assign leaf[327] = f[578] && !f[712] && !f[176] && f[651]; // c3t203i20
	assign leaf[328] = f[578] && !f[712] && f[176] && !f[314]; // c3t203i20
	assign leaf[329] = f[578] && !f[712] && f[176] && f[314]; // c3t203i20
	assign leaf[330] = f[578] && f[712] && !f[461] && !f[372]; // c3t203i20
	assign leaf[331] = f[578] && f[712] && !f[461] && f[372]; // c3t203i20
	assign leaf[332] = f[578] && f[712] && f[461] && !f[206]; // c3t203i20
	assign leaf[333] = f[578] && f[712] && f[461] && f[206]; // c3t203i20
	assign leaf[334] = !f[429] && !f[537] && !f[544] && !f[240]; // c3t213i21
	assign leaf[335] = !f[429] && !f[537] && !f[544] && f[240]; // c3t213i21
	assign leaf[336] = !f[429] && !f[537] && f[544] && !f[489]; // c3t213i21
	assign leaf[337] = !f[429] && !f[537] && f[544] && f[489]; // c3t213i21
	assign leaf[338] = !f[429] && f[537] && !f[326] && !f[382]; // c3t213i21
	assign leaf[339] = !f[429] && f[537] && !f[326] && f[382]; // c3t213i21
	assign leaf[340] = !f[429] && f[537] && f[326] && !f[545]; // c3t213i21
	assign leaf[341] = !f[429] && f[537] && f[326] && f[545]; // c3t213i21
	assign leaf[342] = f[429] && !f[512] && !f[404] && !f[582]; // c3t213i21
	assign leaf[343] = f[429] && !f[512] && !f[404] && f[582]; // c3t213i21
	assign leaf[344] = f[429] && !f[512] && f[404] && !f[370]; // c3t213i21
	assign leaf[345] = f[429] && !f[512] && f[404] && f[370]; // c3t213i21
	assign leaf[346] = f[429] && f[512] && !f[425] && !f[484]; // c3t213i21
	assign leaf[347] = f[429] && f[512] && !f[425] && f[484]; // c3t213i21
	assign leaf[348] = f[429] && f[512] && f[425]; // c3t213i21
	assign leaf[349] = !f[373] && !f[320] && !f[406] && !f[323]; // c3t223i22
	assign leaf[350] = !f[373] && !f[320] && !f[406] && f[323]; // c3t223i22
	assign leaf[351] = !f[373] && !f[320] && f[406] && !f[353]; // c3t223i22
	assign leaf[352] = !f[373] && !f[320] && f[406] && f[353]; // c3t223i22
	assign leaf[353] = !f[373] && f[320] && !f[294] && !f[174]; // c3t223i22
	assign leaf[354] = !f[373] && f[320] && !f[294] && f[174]; // c3t223i22
	assign leaf[355] = !f[373] && f[320] && f[294] && !f[431]; // c3t223i22
	assign leaf[356] = !f[373] && f[320] && f[294] && f[431]; // c3t223i22
	assign leaf[357] = f[373] && !f[321] && !f[200] && !f[345]; // c3t223i22
	assign leaf[358] = f[373] && !f[321] && !f[200] && f[345]; // c3t223i22
	assign leaf[359] = f[373] && !f[321] && f[200] && !f[240]; // c3t223i22
	assign leaf[360] = f[373] && !f[321] && f[200] && f[240]; // c3t223i22
	assign leaf[361] = f[373] && f[321] && !f[327] && !f[246]; // c3t223i22
	assign leaf[362] = f[373] && f[321] && !f[327] && f[246]; // c3t223i22
	assign leaf[363] = f[373] && f[321] && f[327] && !f[455]; // c3t223i22
	assign leaf[364] = f[373] && f[321] && f[327] && f[455]; // c3t223i22
	assign leaf[365] = !f[386] && !f[485] && !f[654] && !f[569]; // c3t233i23
	assign leaf[366] = !f[386] && !f[485] && !f[654] && f[569]; // c3t233i23
	assign leaf[367] = !f[386] && !f[485] && f[654] && !f[543]; // c3t233i23
	assign leaf[368] = !f[386] && !f[485] && f[654] && f[543]; // c3t233i23
	assign leaf[369] = !f[386] && f[485] && !f[480] && !f[710]; // c3t233i23
	assign leaf[370] = !f[386] && f[485] && !f[480] && f[710]; // c3t233i23
	assign leaf[371] = !f[386] && f[485] && f[480] && !f[570]; // c3t233i23
	assign leaf[372] = !f[386] && f[485] && f[480] && f[570]; // c3t233i23
	assign leaf[373] = f[386] && !f[355]; // c3t233i23
	assign leaf[374] = f[386] && f[355] && !f[294] && !f[564]; // c3t233i23
	assign leaf[375] = f[386] && f[355] && !f[294] && f[564]; // c3t233i23
	assign leaf[376] = f[386] && f[355] && f[294] && !f[150]; // c3t233i23
	assign leaf[377] = f[386] && f[355] && f[294] && f[150]; // c3t233i23
	assign leaf[378] = !f[357] && !f[123] && !f[682] && !f[202]; // c3t243i24
	assign leaf[379] = !f[357] && !f[123] && !f[682] && f[202]; // c3t243i24
	assign leaf[380] = !f[357] && !f[123] && f[682] && !f[572]; // c3t243i24
	assign leaf[381] = !f[357] && !f[123] && f[682] && f[572]; // c3t243i24
	assign leaf[382] = !f[357] && f[123] && !f[234] && !f[260]; // c3t243i24
	assign leaf[383] = !f[357] && f[123] && !f[234] && f[260]; // c3t243i24
	assign leaf[384] = !f[357] && f[123] && f[234] && !f[147]; // c3t243i24
	assign leaf[385] = !f[357] && f[123] && f[234] && f[147]; // c3t243i24
	assign leaf[386] = f[357] && !f[355] && !f[488]; // c3t243i24
	assign leaf[387] = f[357] && !f[355] && f[488] && !f[213]; // c3t243i24
	assign leaf[388] = f[357] && !f[355] && f[488] && f[213]; // c3t243i24
	assign leaf[389] = f[357] && f[355] && !f[399] && !f[239]; // c3t243i24
	assign leaf[390] = f[357] && f[355] && !f[399] && f[239]; // c3t243i24
	assign leaf[391] = f[357] && f[355] && f[399] && !f[160]; // c3t243i24
	assign leaf[392] = f[357] && f[355] && f[399] && f[160]; // c3t243i24
	assign leaf[393] = !f[429] && !f[124] && !f[406] && !f[465]; // c3t253i25
	assign leaf[394] = !f[429] && !f[124] && !f[406] && f[465]; // c3t253i25
	assign leaf[395] = !f[429] && !f[124] && f[406] && !f[347]; // c3t253i25
	assign leaf[396] = !f[429] && !f[124] && f[406] && f[347]; // c3t253i25
	assign leaf[397] = !f[429] && f[124] && !f[207] && !f[233]; // c3t253i25
	assign leaf[398] = !f[429] && f[124] && !f[207] && f[233]; // c3t253i25
	assign leaf[399] = !f[429] && f[124] && f[207] && !f[210]; // c3t253i25
	assign leaf[400] = !f[429] && f[124] && f[207] && f[210]; // c3t253i25
	assign leaf[401] = f[429] && !f[511] && !f[404] && !f[554]; // c3t253i25
	assign leaf[402] = f[429] && !f[511] && !f[404] && f[554]; // c3t253i25
	assign leaf[403] = f[429] && !f[511] && f[404] && !f[344]; // c3t253i25
	assign leaf[404] = f[429] && !f[511] && f[404] && f[344]; // c3t253i25
	assign leaf[405] = f[429] && f[511] && !f[425] && !f[456]; // c3t253i25
	assign leaf[406] = f[429] && f[511] && !f[425] && f[456]; // c3t253i25
	assign leaf[407] = f[429] && f[511] && f[425] && !f[572]; // c3t253i25
	assign leaf[408] = f[429] && f[511] && f[425] && f[572]; // c3t253i25
	assign leaf[409] = !f[712] && !f[120] && !f[242] && !f[239]; // c3t263i26
	assign leaf[410] = !f[712] && !f[120] && !f[242] && f[239]; // c3t263i26
	assign leaf[411] = !f[712] && !f[120] && f[242] && !f[157]; // c3t263i26
	assign leaf[412] = !f[712] && !f[120] && f[242] && f[157]; // c3t263i26
	assign leaf[413] = !f[712] && f[120] && !f[632] && !f[293]; // c3t263i26
	assign leaf[414] = !f[712] && f[120] && !f[632] && f[293]; // c3t263i26
	assign leaf[415] = !f[712] && f[120] && f[632] && !f[235]; // c3t263i26
	assign leaf[416] = !f[712] && f[120] && f[632] && f[235]; // c3t263i26
	assign leaf[417] = f[712] && !f[601] && !f[376] && !f[435]; // c3t263i26
	assign leaf[418] = f[712] && !f[601] && !f[376] && f[435]; // c3t263i26
	assign leaf[419] = f[712] && !f[601] && f[376] && !f[232]; // c3t263i26
	assign leaf[420] = f[712] && !f[601] && f[376] && f[232]; // c3t263i26
	assign leaf[421] = f[712] && f[601] && !f[659] && !f[738]; // c3t263i26
	assign leaf[422] = f[712] && f[601] && !f[659] && f[738]; // c3t263i26
	assign leaf[423] = f[712] && f[601] && f[659] && !f[374]; // c3t263i26
	assign leaf[424] = f[712] && f[601] && f[659] && f[374]; // c3t263i26
	assign leaf[425] = !f[200] && !f[373] && !f[320] && !f[681]; // c3t273i27
	assign leaf[426] = !f[200] && !f[373] && !f[320] && f[681]; // c3t273i27
	assign leaf[427] = !f[200] && !f[373] && f[320] && !f[267]; // c3t273i27
	assign leaf[428] = !f[200] && !f[373] && f[320] && f[267]; // c3t273i27
	assign leaf[429] = !f[200] && f[373] && !f[321] && !f[345]; // c3t273i27
	assign leaf[430] = !f[200] && f[373] && !f[321] && f[345]; // c3t273i27
	assign leaf[431] = !f[200] && f[373] && f[321] && !f[256]; // c3t273i27
	assign leaf[432] = !f[200] && f[373] && f[321] && f[256]; // c3t273i27
	assign leaf[433] = f[200] && !f[314] && !f[298] && !f[410]; // c3t273i27
	assign leaf[434] = f[200] && !f[314] && !f[298] && f[410]; // c3t273i27
	assign leaf[435] = f[200] && !f[314] && f[298] && !f[547]; // c3t273i27
	assign leaf[436] = f[200] && !f[314] && f[298] && f[547]; // c3t273i27
	assign leaf[437] = f[200] && f[314]; // c3t273i27
	assign leaf[438] = !f[429] && !f[98] && !f[467] && !f[571]; // c3t283i28
	assign leaf[439] = !f[429] && !f[98] && !f[467] && f[571]; // c3t283i28
	assign leaf[440] = !f[429] && !f[98] && f[467] && !f[407]; // c3t283i28
	assign leaf[441] = !f[429] && !f[98] && f[467] && f[407]; // c3t283i28
	assign leaf[442] = !f[429] && f[98] && !f[208] && !f[431]; // c3t283i28
	assign leaf[443] = !f[429] && f[98] && !f[208] && f[431]; // c3t283i28
	assign leaf[444] = !f[429] && f[98] && f[208] && !f[297]; // c3t283i28
	assign leaf[445] = !f[429] && f[98] && f[208] && f[297]; // c3t283i28
	assign leaf[446] = f[429] && !f[512] && !f[482] && !f[344]; // c3t283i28
	assign leaf[447] = f[429] && !f[512] && !f[482] && f[344]; // c3t283i28
	assign leaf[448] = f[429] && !f[512] && f[482] && !f[686]; // c3t283i28
	assign leaf[449] = f[429] && !f[512] && f[482] && f[686]; // c3t283i28
	assign leaf[450] = f[429] && f[512] && !f[453] && !f[201]; // c3t283i28
	assign leaf[451] = f[429] && f[512] && !f[453] && f[201]; // c3t283i28
	assign leaf[452] = f[429] && f[512] && f[453] && !f[432]; // c3t283i28
	assign leaf[453] = f[429] && f[512] && f[453] && f[432]; // c3t283i28
	assign leaf[454] = !f[678] && !f[147] && !f[318] && !f[292]; // c3t293i29
	assign leaf[455] = !f[678] && !f[147] && !f[318] && f[292]; // c3t293i29
	assign leaf[456] = !f[678] && !f[147] && f[318] && !f[293]; // c3t293i29
	assign leaf[457] = !f[678] && !f[147] && f[318] && f[293]; // c3t293i29
	assign leaf[458] = !f[678] && f[147] && !f[633] && !f[319]; // c3t293i29
	assign leaf[459] = !f[678] && f[147] && !f[633] && f[319]; // c3t293i29
	assign leaf[460] = !f[678] && f[147] && f[633] && !f[314]; // c3t293i29
	assign leaf[461] = !f[678] && f[147] && f[633] && f[314]; // c3t293i29
	assign leaf[462] = f[678] && !f[568] && !f[460] && !f[323]; // c3t293i29
	assign leaf[463] = f[678] && !f[568] && !f[460] && f[323]; // c3t293i29
	assign leaf[464] = f[678] && !f[568] && f[460] && !f[538]; // c3t293i29
	assign leaf[465] = f[678] && !f[568] && f[460] && f[538]; // c3t293i29
	assign leaf[466] = f[678] && f[568] && !f[514]; // c3t293i29
	assign leaf[467] = f[678] && f[568] && f[514]; // c3t293i29
	assign leaf[468] = !f[429] && !f[549] && !f[487] && !f[553]; // c3t303i30
	assign leaf[469] = !f[429] && !f[549] && !f[487] && f[553]; // c3t303i30
	assign leaf[470] = !f[429] && !f[549] && f[487] && !f[716]; // c3t303i30
	assign leaf[471] = !f[429] && !f[549] && f[487] && f[716]; // c3t303i30
	assign leaf[472] = !f[429] && f[549] && !f[712] && !f[263]; // c3t303i30
	assign leaf[473] = !f[429] && f[549] && !f[712] && f[263]; // c3t303i30
	assign leaf[474] = !f[429] && f[549] && f[712] && !f[320]; // c3t303i30
	assign leaf[475] = !f[429] && f[549] && f[712] && f[320]; // c3t303i30
	assign leaf[476] = f[429] && !f[433] && !f[516] && !f[482]; // c3t303i30
	assign leaf[477] = f[429] && !f[433] && !f[516] && f[482]; // c3t303i30
	assign leaf[478] = f[429] && !f[433] && f[516] && !f[464]; // c3t303i30
	assign leaf[479] = f[429] && !f[433] && f[516] && f[464]; // c3t303i30
	assign leaf[480] = f[429] && f[433] && !f[580] && !f[549]; // c3t303i30
	assign leaf[481] = f[429] && f[433] && !f[580] && f[549]; // c3t303i30
	assign leaf[482] = f[429] && f[433] && f[580] && !f[370]; // c3t303i30
	assign leaf[483] = f[429] && f[433] && f[580] && f[370]; // c3t303i30
	assign leaf[484] = !f[399] && !f[536] && !f[551] && !f[125]; // c3t313i31
	assign leaf[485] = !f[399] && !f[536] && !f[551] && f[125]; // c3t313i31
	assign leaf[486] = !f[399] && !f[536] && f[551] && !f[238]; // c3t313i31
	assign leaf[487] = !f[399] && !f[536] && f[551] && f[238]; // c3t313i31
	assign leaf[488] = !f[399] && f[536] && !f[299] && !f[376]; // c3t313i31
	assign leaf[489] = !f[399] && f[536] && !f[299] && f[376]; // c3t313i31
	assign leaf[490] = !f[399] && f[536] && f[299] && !f[483]; // c3t313i31
	assign leaf[491] = !f[399] && f[536] && f[299] && f[483]; // c3t313i31
	assign leaf[492] = f[399] && !f[294] && !f[412] && !f[288]; // c3t313i31
	assign leaf[493] = f[399] && !f[294] && !f[412] && f[288]; // c3t313i31
	assign leaf[494] = f[399] && !f[294] && f[412] && !f[296]; // c3t313i31
	assign leaf[495] = f[399] && !f[294] && f[412] && f[296]; // c3t313i31
	assign leaf[496] = f[399] && f[294] && !f[288] && !f[526]; // c3t313i31
	assign leaf[497] = f[399] && f[294] && !f[288] && f[526]; // c3t313i31
	assign leaf[498] = f[399] && f[294] && f[288] && !f[516]; // c3t313i31
	assign leaf[499] = f[399] && f[294] && f[288] && f[516]; // c3t313i31
	assign leaf[500] = !f[370] && !f[346] && !f[320] && !f[372]; // c3t323i32
	assign leaf[501] = !f[370] && !f[346] && !f[320] && f[372]; // c3t323i32
	assign leaf[502] = !f[370] && !f[346] && f[320] && !f[292]; // c3t323i32
	assign leaf[503] = !f[370] && !f[346] && f[320] && f[292]; // c3t323i32
	assign leaf[504] = !f[370] && f[346] && !f[321] && !f[375]; // c3t323i32
	assign leaf[505] = !f[370] && f[346] && !f[321] && f[375]; // c3t323i32
	assign leaf[506] = !f[370] && f[346] && f[321] && !f[263]; // c3t323i32
	assign leaf[507] = !f[370] && f[346] && f[321] && f[263]; // c3t323i32
	assign leaf[508] = f[370] && !f[711] && !f[314] && !f[377]; // c3t323i32
	assign leaf[509] = f[370] && !f[711] && !f[314] && f[377]; // c3t323i32
	assign leaf[510] = f[370] && !f[711] && f[314] && !f[284]; // c3t323i32
	assign leaf[511] = f[370] && !f[711] && f[314] && f[284]; // c3t323i32
	assign leaf[512] = f[370] && f[711]; // c3t323i32
	assign leaf[513] = !f[712] && !f[535] && !f[657] && !f[458]; // c3t333i33
	assign leaf[514] = !f[712] && !f[535] && !f[657] && f[458]; // c3t333i33
	assign leaf[515] = !f[712] && !f[535] && f[657] && !f[709]; // c3t333i33
	assign leaf[516] = !f[712] && !f[535] && f[657] && f[709]; // c3t333i33
	assign leaf[517] = !f[712] && f[535] && !f[458] && !f[441]; // c3t333i33
	assign leaf[518] = !f[712] && f[535] && !f[458] && f[441]; // c3t333i33
	assign leaf[519] = !f[712] && f[535] && f[458] && !f[510]; // c3t333i33
	assign leaf[520] = !f[712] && f[535] && f[458] && f[510]; // c3t333i33
	assign leaf[521] = f[712] && !f[573] && !f[489] && !f[343]; // c3t333i33
	assign leaf[522] = f[712] && !f[573] && !f[489] && f[343]; // c3t333i33
	assign leaf[523] = f[712] && !f[573] && f[489] && !f[598]; // c3t333i33
	assign leaf[524] = f[712] && !f[573] && f[489] && f[598]; // c3t333i33
	assign leaf[525] = f[712] && f[573] && !f[488] && !f[429]; // c3t333i33
	assign leaf[526] = f[712] && f[573] && !f[488] && f[429]; // c3t333i33
	assign leaf[527] = f[712] && f[573] && f[488] && !f[599]; // c3t333i33
	assign leaf[528] = f[712] && f[573] && f[488] && f[599]; // c3t333i33
	assign leaf[529] = !f[712] && !f[649] && !f[173] && !f[480]; // c3t343i34
	assign leaf[530] = !f[712] && !f[649] && !f[173] && f[480]; // c3t343i34
	assign leaf[531] = !f[712] && !f[649] && f[173] && !f[553]; // c3t343i34
	assign leaf[532] = !f[712] && !f[649] && f[173] && f[553]; // c3t343i34
	assign leaf[533] = !f[712] && f[649] && !f[539] && !f[320]; // c3t343i34
	assign leaf[534] = !f[712] && f[649] && !f[539] && f[320]; // c3t343i34
	assign leaf[535] = !f[712] && f[649] && f[539] && !f[375]; // c3t343i34
	assign leaf[536] = !f[712] && f[649] && f[539] && f[375]; // c3t343i34
	assign leaf[537] = f[712] && !f[600] && !f[489] && !f[519]; // c3t343i34
	assign leaf[538] = f[712] && !f[600] && !f[489] && f[519]; // c3t343i34
	assign leaf[539] = f[712] && !f[600] && f[489] && !f[403]; // c3t343i34
	assign leaf[540] = f[712] && !f[600] && f[489] && f[403]; // c3t343i34
	assign leaf[541] = f[712] && f[600] && !f[287] && !f[328]; // c3t343i34
	assign leaf[542] = f[712] && f[600] && !f[287] && f[328]; // c3t343i34
	assign leaf[543] = f[712] && f[600] && f[287]; // c3t343i34
	assign leaf[544] = !f[373] && !f[523] && !f[320] && !f[327]; // c3t353i35
	assign leaf[545] = !f[373] && !f[523] && !f[320] && f[327]; // c3t353i35
	assign leaf[546] = !f[373] && !f[523] && f[320] && !f[126]; // c3t353i35
	assign leaf[547] = !f[373] && !f[523] && f[320] && f[126]; // c3t353i35
	assign leaf[548] = !f[373] && f[523] && !f[238] && !f[263]; // c3t353i35
	assign leaf[549] = !f[373] && f[523] && !f[238] && f[263]; // c3t353i35
	assign leaf[550] = !f[373] && f[523] && f[238] && !f[161]; // c3t353i35
	assign leaf[551] = !f[373] && f[523] && f[238] && f[161]; // c3t353i35
	assign leaf[552] = f[373] && !f[288] && !f[526] && !f[154]; // c3t353i35
	assign leaf[553] = f[373] && !f[288] && !f[526] && f[154]; // c3t353i35
	assign leaf[554] = f[373] && !f[288] && f[526] && !f[293]; // c3t353i35
	assign leaf[555] = f[373] && !f[288] && f[526] && f[293]; // c3t353i35
	assign leaf[556] = f[373] && f[288] && !f[264] && !f[316]; // c3t353i35
	assign leaf[557] = f[373] && f[288] && !f[264] && f[316]; // c3t353i35
	assign leaf[558] = f[373] && f[288] && f[264] && !f[469]; // c3t353i35
	assign leaf[559] = f[373] && f[288] && f[264] && f[469]; // c3t353i35
	assign leaf[560] = !f[386] && !f[269] && !f[129] && !f[491]; // c3t363i36
	assign leaf[561] = !f[386] && !f[269] && !f[129] && f[491]; // c3t363i36
	assign leaf[562] = !f[386] && !f[269] && f[129] && !f[272]; // c3t363i36
	assign leaf[563] = !f[386] && !f[269] && f[129] && f[272]; // c3t363i36
	assign leaf[564] = !f[386] && f[269] && !f[99] && !f[572]; // c3t363i36
	assign leaf[565] = !f[386] && f[269] && !f[99] && f[572]; // c3t363i36
	assign leaf[566] = !f[386] && f[269] && f[99] && !f[179]; // c3t363i36
	assign leaf[567] = !f[386] && f[269] && f[99] && f[179]; // c3t363i36
	assign leaf[568] = f[386] && !f[354]; // c3t363i36
	assign leaf[569] = f[386] && f[354] && !f[149] && !f[381]; // c3t363i36
	assign leaf[570] = f[386] && f[354] && !f[149] && f[381]; // c3t363i36
	assign leaf[571] = f[386] && f[354] && f[149] && !f[267]; // c3t363i36
	assign leaf[572] = f[386] && f[354] && f[149] && f[267]; // c3t363i36
	assign leaf[573] = !f[708] && !f[550] && !f[553] && !f[98]; // c3t373i37
	assign leaf[574] = !f[708] && !f[550] && !f[553] && f[98]; // c3t373i37
	assign leaf[575] = !f[708] && !f[550] && f[553] && !f[547]; // c3t373i37
	assign leaf[576] = !f[708] && !f[550] && f[553] && f[547]; // c3t373i37
	assign leaf[577] = !f[708] && f[550] && !f[401] && !f[544]; // c3t373i37
	assign leaf[578] = !f[708] && f[550] && !f[401] && f[544]; // c3t373i37
	assign leaf[579] = !f[708] && f[550] && f[401] && !f[455]; // c3t373i37
	assign leaf[580] = !f[708] && f[550] && f[401] && f[455]; // c3t373i37
	assign leaf[581] = f[708] && !f[576] && !f[599] && !f[293]; // c3t373i37
	assign leaf[582] = f[708] && !f[576] && !f[599] && f[293]; // c3t373i37
	assign leaf[583] = f[708] && !f[576] && f[599] && !f[516]; // c3t373i37
	assign leaf[584] = f[708] && !f[576] && f[599] && f[516]; // c3t373i37
	assign leaf[585] = f[708] && f[576] && !f[376]; // c3t373i37
	assign leaf[586] = f[708] && f[576] && f[376] && !f[380]; // c3t373i37
	assign leaf[587] = f[708] && f[576] && f[376] && f[380]; // c3t373i37
	assign leaf[588] = !f[457] && !f[96] && !f[406] && !f[461]; // c3t383i38
	assign leaf[589] = !f[457] && !f[96] && !f[406] && f[461]; // c3t383i38
	assign leaf[590] = !f[457] && !f[96] && f[406] && !f[300]; // c3t383i38
	assign leaf[591] = !f[457] && !f[96] && f[406] && f[300]; // c3t383i38
	assign leaf[592] = !f[457] && f[96] && !f[265] && !f[568]; // c3t383i38
	assign leaf[593] = !f[457] && f[96] && !f[265] && f[568]; // c3t383i38
	assign leaf[594] = !f[457] && f[96] && f[265] && !f[180]; // c3t383i38
	assign leaf[595] = !f[457] && f[96] && f[265] && f[180]; // c3t383i38
	assign leaf[596] = f[457] && !f[235] && !f[578] && !f[508]; // c3t383i38
	assign leaf[597] = f[457] && !f[235] && !f[578] && f[508]; // c3t383i38
	assign leaf[598] = f[457] && !f[235] && f[578] && !f[324]; // c3t383i38
	assign leaf[599] = f[457] && !f[235] && f[578] && f[324]; // c3t383i38
	assign leaf[600] = f[457] && f[235] && !f[406] && !f[598]; // c3t383i38
	assign leaf[601] = f[457] && f[235] && !f[406] && f[598]; // c3t383i38
	assign leaf[602] = f[457] && f[235] && f[406] && !f[346]; // c3t383i38
	assign leaf[603] = f[457] && f[235] && f[406] && f[346]; // c3t383i38
	assign leaf[604] = !f[358] && !f[486] && !f[456] && !f[595]; // c3t393i39
	assign leaf[605] = !f[358] && !f[486] && !f[456] && f[595]; // c3t393i39
	assign leaf[606] = !f[358] && !f[486] && f[456] && !f[299]; // c3t393i39
	assign leaf[607] = !f[358] && !f[486] && f[456] && f[299]; // c3t393i39
	assign leaf[608] = !f[358] && f[486] && !f[716] && !f[577]; // c3t393i39
	assign leaf[609] = !f[358] && f[486] && !f[716] && f[577]; // c3t393i39
	assign leaf[610] = !f[358] && f[486] && f[716] && !f[438]; // c3t393i39
	assign leaf[611] = !f[358] && f[486] && f[716] && f[438]; // c3t393i39
	assign leaf[612] = f[358] && !f[291] && !f[650]; // c3t393i39
	assign leaf[613] = f[358] && !f[291] && f[650]; // c3t393i39
	assign leaf[614] = f[358] && f[291] && !f[582] && !f[319]; // c3t393i39
	assign leaf[615] = f[358] && f[291] && !f[582] && f[319]; // c3t393i39
	assign leaf[616] = f[358] && f[291] && f[582]; // c3t393i39
	assign leaf[617] = !f[210] && !f[234] && !f[156] && !f[525]; // c3t403i40
	assign leaf[618] = !f[210] && !f[234] && !f[156] && f[525]; // c3t403i40
	assign leaf[619] = !f[210] && !f[234] && f[156] && !f[236]; // c3t403i40
	assign leaf[620] = !f[210] && !f[234] && f[156] && f[236]; // c3t403i40
	assign leaf[621] = !f[210] && f[234] && !f[151] && !f[491]; // c3t403i40
	assign leaf[622] = !f[210] && f[234] && !f[151] && f[491]; // c3t403i40
	assign leaf[623] = !f[210] && f[234] && f[151] && !f[258]; // c3t403i40
	assign leaf[624] = !f[210] && f[234] && f[151] && f[258]; // c3t403i40
	assign leaf[625] = f[210] && !f[346] && !f[572] && !f[489]; // c3t403i40
	assign leaf[626] = f[210] && !f[346] && !f[572] && f[489]; // c3t403i40
	assign leaf[627] = f[210] && !f[346] && f[572] && !f[536]; // c3t403i40
	assign leaf[628] = f[210] && !f[346] && f[572] && f[536]; // c3t403i40
	assign leaf[629] = f[210] && f[346] && !f[442] && !f[375]; // c3t403i40
	assign leaf[630] = f[210] && f[346] && !f[442] && f[375]; // c3t403i40
	assign leaf[631] = f[210] && f[346] && f[442] && !f[314]; // c3t403i40
	assign leaf[632] = f[210] && f[346] && f[442] && f[314]; // c3t403i40
	assign leaf[633] = !f[269] && !f[513] && !f[497] && !f[299]; // c3t413i41
	assign leaf[634] = !f[269] && !f[513] && !f[497] && f[299]; // c3t413i41
	assign leaf[635] = !f[269] && !f[513] && f[497] && !f[265]; // c3t413i41
	assign leaf[636] = !f[269] && !f[513] && f[497] && f[265]; // c3t413i41
	assign leaf[637] = !f[269] && f[513] && !f[509] && !f[523]; // c3t413i41
	assign leaf[638] = !f[269] && f[513] && !f[509] && f[523]; // c3t413i41
	assign leaf[639] = !f[269] && f[513] && f[509] && !f[462]; // c3t413i41
	assign leaf[640] = !f[269] && f[513] && f[509] && f[462]; // c3t413i41
	assign leaf[641] = f[269] && !f[341] && !f[323] && !f[433]; // c3t413i41
	assign leaf[642] = f[269] && !f[341] && !f[323] && f[433]; // c3t413i41
	assign leaf[643] = f[269] && !f[341] && f[323] && !f[494]; // c3t413i41
	assign leaf[644] = f[269] && !f[341] && f[323] && f[494]; // c3t413i41
	assign leaf[645] = f[269] && f[341] && !f[656]; // c3t413i41
	assign leaf[646] = f[269] && f[341] && f[656] && !f[399]; // c3t413i41
	assign leaf[647] = f[269] && f[341] && f[656] && f[399]; // c3t413i41
	assign leaf[648] = !f[371] && !f[211] && !f[235] && !f[156]; // c3t423i42
	assign leaf[649] = !f[371] && !f[211] && !f[235] && f[156]; // c3t423i42
	assign leaf[650] = !f[371] && !f[211] && f[235] && !f[202]; // c3t423i42
	assign leaf[651] = !f[371] && !f[211] && f[235] && f[202]; // c3t423i42
	assign leaf[652] = !f[371] && f[211] && !f[131] && !f[549]; // c3t423i42
	assign leaf[653] = !f[371] && f[211] && !f[131] && f[549]; // c3t423i42
	assign leaf[654] = !f[371] && f[211] && f[131] && !f[266]; // c3t423i42
	assign leaf[655] = !f[371] && f[211] && f[131] && f[266]; // c3t423i42
	assign leaf[656] = f[371] && !f[315] && !f[313] && !f[481]; // c3t423i42
	assign leaf[657] = f[371] && !f[315] && !f[313] && f[481]; // c3t423i42
	assign leaf[658] = f[371] && !f[315] && f[313]; // c3t423i42
	assign leaf[659] = f[371] && f[315] && !f[232] && !f[351]; // c3t423i42
	assign leaf[660] = f[371] && f[315] && !f[232] && f[351]; // c3t423i42
	assign leaf[661] = f[371] && f[315] && f[232] && !f[689]; // c3t423i42
	assign leaf[662] = f[371] && f[315] && f[232] && f[689]; // c3t423i42
	assign leaf[663] = !f[708] && !f[120] && !f[318] && !f[344]; // c3t433i43
	assign leaf[664] = !f[708] && !f[120] && !f[318] && f[344]; // c3t433i43
	assign leaf[665] = !f[708] && !f[120] && f[318] && !f[293]; // c3t433i43
	assign leaf[666] = !f[708] && !f[120] && f[318] && f[293]; // c3t433i43
	assign leaf[667] = !f[708] && f[120] && !f[292] && !f[345]; // c3t433i43
	assign leaf[668] = !f[708] && f[120] && !f[292] && f[345]; // c3t433i43
	assign leaf[669] = !f[708] && f[120] && f[292] && !f[260]; // c3t433i43
	assign leaf[670] = !f[708] && f[120] && f[292] && f[260]; // c3t433i43
	assign leaf[671] = f[708] && !f[599] && !f[463] && !f[377]; // c3t433i43
	assign leaf[672] = f[708] && !f[599] && !f[463] && f[377]; // c3t433i43
	assign leaf[673] = f[708] && !f[599] && f[463] && !f[382]; // c3t433i43
	assign leaf[674] = f[708] && !f[599] && f[463] && f[382]; // c3t433i43
	assign leaf[675] = f[708] && f[599] && !f[602]; // c3t433i43
	assign leaf[676] = f[708] && f[599] && f[602]; // c3t433i43
	assign leaf[677] = !f[427] && !f[486] && !f[124] && !f[554]; // c3t443i44
	assign leaf[678] = !f[427] && !f[486] && !f[124] && f[554]; // c3t443i44
	assign leaf[679] = !f[427] && !f[486] && f[124] && !f[207]; // c3t443i44
	assign leaf[680] = !f[427] && !f[486] && f[124] && f[207]; // c3t443i44
	assign leaf[681] = !f[427] && f[486] && !f[541] && !f[542]; // c3t443i44
	assign leaf[682] = !f[427] && f[486] && !f[541] && f[542]; // c3t443i44
	assign leaf[683] = !f[427] && f[486] && f[541] && !f[483]; // c3t443i44
	assign leaf[684] = !f[427] && f[486] && f[541] && f[483]; // c3t443i44
	assign leaf[685] = f[427] && !f[158] && !f[710] && !f[466]; // c3t443i44
	assign leaf[686] = f[427] && !f[158] && !f[710] && f[466]; // c3t443i44
	assign leaf[687] = f[427] && !f[158] && f[710]; // c3t443i44
	assign leaf[688] = f[427] && f[158] && !f[356] && !f[494]; // c3t443i44
	assign leaf[689] = f[427] && f[158] && !f[356] && f[494]; // c3t443i44
	assign leaf[690] = f[427] && f[158] && f[356] && !f[486]; // c3t443i44
	assign leaf[691] = f[427] && f[158] && f[356] && f[486]; // c3t443i44
	assign leaf[692] = !f[451] && !f[133] && !f[591] && !f[210]; // c3t453i45
	assign leaf[693] = !f[451] && !f[133] && !f[591] && f[210]; // c3t453i45
	assign leaf[694] = !f[451] && !f[133] && f[591] && !f[404]; // c3t453i45
	assign leaf[695] = !f[451] && !f[133] && f[591] && f[404]; // c3t453i45
	assign leaf[696] = !f[451] && f[133] && !f[272] && !f[179]; // c3t453i45
	assign leaf[697] = !f[451] && f[133] && !f[272] && f[179]; // c3t453i45
	assign leaf[698] = !f[451] && f[133] && f[272] && !f[462]; // c3t453i45
	assign leaf[699] = !f[451] && f[133] && f[272] && f[462]; // c3t453i45
	assign leaf[700] = f[451] && !f[352]; // c3t453i45
	assign leaf[701] = f[451] && f[352] && !f[159]; // c3t453i45
	assign leaf[702] = f[451] && f[352] && f[159]; // c3t453i45
	assign leaf[703] = !f[458] && !f[566] && !f[266] && !f[355]; // c3t463i46
	assign leaf[704] = !f[458] && !f[566] && !f[266] && f[355]; // c3t463i46
	assign leaf[705] = !f[458] && !f[566] && f[266] && !f[468]; // c3t463i46
	assign leaf[706] = !f[458] && !f[566] && f[266] && f[468]; // c3t463i46
	assign leaf[707] = !f[458] && f[566] && !f[517] && !f[455]; // c3t463i46
	assign leaf[708] = !f[458] && f[566] && !f[517] && f[455]; // c3t463i46
	assign leaf[709] = !f[458] && f[566] && f[517] && !f[621]; // c3t463i46
	assign leaf[710] = !f[458] && f[566] && f[517] && f[621]; // c3t463i46
	assign leaf[711] = f[458] && !f[489] && !f[540] && !f[653]; // c3t463i46
	assign leaf[712] = f[458] && !f[489] && !f[540] && f[653]; // c3t463i46
	assign leaf[713] = f[458] && !f[489] && f[540] && !f[372]; // c3t463i46
	assign leaf[714] = f[458] && !f[489] && f[540] && f[372]; // c3t463i46
	assign leaf[715] = f[458] && f[489] && !f[605] && !f[436]; // c3t463i46
	assign leaf[716] = f[458] && f[489] && !f[605] && f[436]; // c3t463i46
	assign leaf[717] = f[458] && f[489] && f[605] && !f[346]; // c3t463i46
	assign leaf[718] = f[458] && f[489] && f[605] && f[346]; // c3t463i46
	assign leaf[719] = !f[712] && !f[377] && !f[537] && !f[571]; // c3t473i47
	assign leaf[720] = !f[712] && !f[377] && !f[537] && f[571]; // c3t473i47
	assign leaf[721] = !f[712] && !f[377] && f[537] && !f[209]; // c3t473i47
	assign leaf[722] = !f[712] && !f[377] && f[537] && f[209]; // c3t473i47
	assign leaf[723] = !f[712] && f[377] && !f[484] && !f[318]; // c3t473i47
	assign leaf[724] = !f[712] && f[377] && !f[484] && f[318]; // c3t473i47
	assign leaf[725] = !f[712] && f[377] && f[484] && !f[515]; // c3t473i47
	assign leaf[726] = !f[712] && f[377] && f[484] && f[515]; // c3t473i47
	assign leaf[727] = f[712] && !f[600] && !f[319] && !f[345]; // c3t473i47
	assign leaf[728] = f[712] && !f[600] && !f[319] && f[345]; // c3t473i47
	assign leaf[729] = f[712] && !f[600] && f[319] && !f[348]; // c3t473i47
	assign leaf[730] = f[712] && !f[600] && f[319] && f[348]; // c3t473i47
	assign leaf[731] = f[712] && f[600] && !f[317]; // c3t473i47
	assign leaf[732] = f[712] && f[600] && f[317]; // c3t473i47
	assign leaf[733] = !f[161] && !f[655] && !f[464] && !f[548]; // c3t483i48
	assign leaf[734] = !f[161] && !f[655] && !f[464] && f[548]; // c3t483i48
	assign leaf[735] = !f[161] && !f[655] && f[464] && !f[547]; // c3t483i48
	assign leaf[736] = !f[161] && !f[655] && f[464] && f[547]; // c3t483i48
	assign leaf[737] = !f[161] && f[655] && !f[630] && !f[544]; // c3t483i48
	assign leaf[738] = !f[161] && f[655] && !f[630] && f[544]; // c3t483i48
	assign leaf[739] = !f[161] && f[655] && f[630] && !f[710]; // c3t483i48
	assign leaf[740] = !f[161] && f[655] && f[630] && f[710]; // c3t483i48
	assign leaf[741] = f[161] && !f[272] && !f[301] && !f[243]; // c3t483i48
	assign leaf[742] = f[161] && !f[272] && !f[301] && f[243]; // c3t483i48
	assign leaf[743] = f[161] && !f[272] && f[301]; // c3t483i48
	assign leaf[744] = f[161] && f[272] && !f[326] && !f[267]; // c3t483i48
	assign leaf[745] = f[161] && f[272] && !f[326] && f[267]; // c3t483i48
	assign leaf[746] = f[161] && f[272] && f[326] && !f[460]; // c3t483i48
	assign leaf[747] = f[161] && f[272] && f[326] && f[460]; // c3t483i48
	assign leaf[748] = !f[228] && !f[406] && !f[96] && !f[436]; // c3t493i49
	assign leaf[749] = !f[228] && !f[406] && !f[96] && f[436]; // c3t493i49
	assign leaf[750] = !f[228] && !f[406] && f[96] && !f[431]; // c3t493i49
	assign leaf[751] = !f[228] && !f[406] && f[96] && f[431]; // c3t493i49
	assign leaf[752] = !f[228] && f[406] && !f[287] && !f[181]; // c3t493i49
	assign leaf[753] = !f[228] && f[406] && !f[287] && f[181]; // c3t493i49
	assign leaf[754] = !f[228] && f[406] && f[287] && !f[262]; // c3t493i49
	assign leaf[755] = !f[228] && f[406] && f[287] && f[262]; // c3t493i49
	assign leaf[756] = f[228] && !f[375] && !f[439] && !f[630]; // c3t493i49
	assign leaf[757] = f[228] && !f[375] && !f[439] && f[630]; // c3t493i49
	assign leaf[758] = f[228] && !f[375] && f[439] && !f[212]; // c3t493i49
	assign leaf[759] = f[228] && !f[375] && f[439] && f[212]; // c3t493i49
	assign leaf[760] = f[228] && f[375] && !f[344] && !f[293]; // c3t493i49
	assign leaf[761] = f[228] && f[375] && !f[344] && f[293]; // c3t493i49
	assign leaf[762] = f[228] && f[375] && f[344]; // c3t493i49
	assign leaf[763] = !f[429] && !f[544] && !f[489] && !f[459]; // c3t503i50
	assign leaf[764] = !f[429] && !f[544] && !f[489] && f[459]; // c3t503i50
	assign leaf[765] = !f[429] && !f[544] && f[489] && !f[460]; // c3t503i50
	assign leaf[766] = !f[429] && !f[544] && f[489] && f[460]; // c3t503i50
	assign leaf[767] = !f[429] && f[544] && !f[538] && !f[572]; // c3t503i50
	assign leaf[768] = !f[429] && f[544] && !f[538] && f[572]; // c3t503i50
	assign leaf[769] = !f[429] && f[544] && f[538] && !f[294]; // c3t503i50
	assign leaf[770] = !f[429] && f[544] && f[538] && f[294]; // c3t503i50
	assign leaf[771] = f[429] && !f[460] && !f[484] && !f[405]; // c3t503i50
	assign leaf[772] = f[429] && !f[460] && !f[484] && f[405]; // c3t503i50
	assign leaf[773] = f[429] && !f[460] && f[484] && !f[402]; // c3t503i50
	assign leaf[774] = f[429] && !f[460] && f[484] && f[402]; // c3t503i50
	assign leaf[775] = f[429] && f[460] && !f[349] && !f[438]; // c3t503i50
	assign leaf[776] = f[429] && f[460] && !f[349] && f[438]; // c3t503i50
	assign leaf[777] = f[429] && f[460] && f[349] && !f[657]; // c3t503i50
	assign leaf[778] = f[429] && f[460] && f[349] && f[657]; // c3t503i50
	assign leaf[779] = !f[373] && !f[316] && !f[718] && !f[689]; // c3t513i51
	assign leaf[780] = !f[373] && !f[316] && !f[718] && f[689]; // c3t513i51
	assign leaf[781] = !f[373] && !f[316] && f[718] && !f[460]; // c3t513i51
	assign leaf[782] = !f[373] && !f[316] && f[718] && f[460]; // c3t513i51
	assign leaf[783] = !f[373] && f[316] && !f[264] && !f[407]; // c3t513i51
	assign leaf[784] = !f[373] && f[316] && !f[264] && f[407]; // c3t513i51
	assign leaf[785] = !f[373] && f[316] && f[264] && !f[398]; // c3t513i51
	assign leaf[786] = !f[373] && f[316] && f[264] && f[398]; // c3t513i51
	assign leaf[787] = f[373] && !f[289] && !f[315] && !f[607]; // c3t513i51
	assign leaf[788] = f[373] && !f[289] && !f[315] && f[607]; // c3t513i51
	assign leaf[789] = f[373] && !f[289] && f[315] && !f[287]; // c3t513i51
	assign leaf[790] = f[373] && !f[289] && f[315] && f[287]; // c3t513i51
	assign leaf[791] = f[373] && f[289] && !f[264] && !f[317]; // c3t513i51
	assign leaf[792] = f[373] && f[289] && !f[264] && f[317]; // c3t513i51
	assign leaf[793] = f[373] && f[289] && f[264] && !f[183]; // c3t513i51
	assign leaf[794] = f[373] && f[289] && f[264] && f[183]; // c3t513i51
	assign leaf[795] = !f[401] && !f[716] && !f[459] && !f[537]; // c3t523i52
	assign leaf[796] = !f[401] && !f[716] && !f[459] && f[537]; // c3t523i52
	assign leaf[797] = !f[401] && !f[716] && f[459] && !f[570]; // c3t523i52
	assign leaf[798] = !f[401] && !f[716] && f[459] && f[570]; // c3t523i52
	assign leaf[799] = !f[401] && f[716] && !f[433] && !f[576]; // c3t523i52
	assign leaf[800] = !f[401] && f[716] && !f[433] && f[576]; // c3t523i52
	assign leaf[801] = !f[401] && f[716] && f[433] && !f[347]; // c3t523i52
	assign leaf[802] = !f[401] && f[716] && f[433] && f[347]; // c3t523i52
	assign leaf[803] = f[401] && !f[482] && !f[344] && !f[513]; // c3t523i52
	assign leaf[804] = f[401] && !f[482] && !f[344] && f[513]; // c3t523i52
	assign leaf[805] = f[401] && !f[482] && f[344] && !f[347]; // c3t523i52
	assign leaf[806] = f[401] && !f[482] && f[344] && f[347]; // c3t523i52
	assign leaf[807] = f[401] && f[482] && !f[538] && !f[578]; // c3t523i52
	assign leaf[808] = f[401] && f[482] && !f[538] && f[578]; // c3t523i52
	assign leaf[809] = f[401] && f[482] && f[538] && !f[541]; // c3t523i52
	assign leaf[810] = f[401] && f[482] && f[538] && f[541]; // c3t523i52
	assign leaf[811] = !f[708] && !f[386] && !f[269] && !f[239]; // c3t533i53
	assign leaf[812] = !f[708] && !f[386] && !f[269] && f[239]; // c3t533i53
	assign leaf[813] = !f[708] && !f[386] && f[269] && !f[101]; // c3t533i53
	assign leaf[814] = !f[708] && !f[386] && f[269] && f[101]; // c3t533i53
	assign leaf[815] = !f[708] && f[386] && !f[355]; // c3t533i53
	assign leaf[816] = !f[708] && f[386] && f[355] && !f[259]; // c3t533i53
	assign leaf[817] = !f[708] && f[386] && f[355] && f[259]; // c3t533i53
	assign leaf[818] = f[708] && !f[599] && !f[274] && !f[488]; // c3t533i53
	assign leaf[819] = f[708] && !f[599] && !f[274] && f[488]; // c3t533i53
	assign leaf[820] = f[708] && !f[599] && f[274]; // c3t533i53
	assign leaf[821] = f[708] && f[599] && !f[602]; // c3t533i53
	assign leaf[822] = f[708] && f[599] && f[602]; // c3t533i53
	assign leaf[823] = !f[712] && !f[370] && !f[480] && !f[678]; // c3t543i54
	assign leaf[824] = !f[712] && !f[370] && !f[480] && f[678]; // c3t543i54
	assign leaf[825] = !f[712] && !f[370] && f[480] && !f[545]; // c3t543i54
	assign leaf[826] = !f[712] && !f[370] && f[480] && f[545]; // c3t543i54
	assign leaf[827] = !f[712] && f[370] && !f[286] && !f[492]; // c3t543i54
	assign leaf[828] = !f[712] && f[370] && !f[286] && f[492]; // c3t543i54
	assign leaf[829] = !f[712] && f[370] && f[286] && !f[316]; // c3t543i54
	assign leaf[830] = !f[712] && f[370] && f[286] && f[316]; // c3t543i54
	assign leaf[831] = f[712] && !f[231] && !f[295] && !f[689]; // c3t543i54
	assign leaf[832] = f[712] && !f[231] && !f[295] && f[689]; // c3t543i54
	assign leaf[833] = f[712] && !f[231] && f[295] && !f[180]; // c3t543i54
	assign leaf[834] = f[712] && !f[231] && f[295] && f[180]; // c3t543i54
	assign leaf[835] = f[712] && f[231] && !f[465] && !f[604]; // c3t543i54
	assign leaf[836] = f[712] && f[231] && !f[465] && f[604]; // c3t543i54
	assign leaf[837] = f[712] && f[231] && f[465] && !f[578]; // c3t543i54
	assign leaf[838] = f[712] && f[231] && f[465] && f[578]; // c3t543i54
	assign leaf[839] = !f[241] && !f[203] && !f[147] && !f[244]; // c3t553i55
	assign leaf[840] = !f[241] && !f[203] && !f[147] && f[244]; // c3t553i55
	assign leaf[841] = !f[241] && !f[203] && f[147] && !f[264]; // c3t553i55
	assign leaf[842] = !f[241] && !f[203] && f[147] && f[264]; // c3t553i55
	assign leaf[843] = !f[241] && f[203] && !f[259] && !f[492]; // c3t553i55
	assign leaf[844] = !f[241] && f[203] && !f[259] && f[492]; // c3t553i55
	assign leaf[845] = !f[241] && f[203] && f[259] && !f[434]; // c3t553i55
	assign leaf[846] = !f[241] && f[203] && f[259] && f[434]; // c3t553i55
	assign leaf[847] = f[241] && !f[347] && !f[290] && !f[372]; // c3t553i55
	assign leaf[848] = f[241] && !f[347] && !f[290] && f[372]; // c3t553i55
	assign leaf[849] = f[241] && !f[347] && f[290] && !f[179]; // c3t553i55
	assign leaf[850] = f[241] && !f[347] && f[290] && f[179]; // c3t553i55
	assign leaf[851] = f[241] && f[347] && !f[264] && !f[289]; // c3t553i55
	assign leaf[852] = f[241] && f[347] && !f[264] && f[289]; // c3t553i55
	assign leaf[853] = f[241] && f[347] && f[264] && !f[295]; // c3t553i55
	assign leaf[854] = f[241] && f[347] && f[264] && f[295]; // c3t553i55
	assign leaf[855] = !f[369] && !f[402] && !f[544] && !f[211]; // c3t563i56
	assign leaf[856] = !f[369] && !f[402] && !f[544] && f[211]; // c3t563i56
	assign leaf[857] = !f[369] && !f[402] && f[544] && !f[547]; // c3t563i56
	assign leaf[858] = !f[369] && !f[402] && f[544] && f[547]; // c3t563i56
	assign leaf[859] = !f[369] && f[402] && !f[526] && !f[318]; // c3t563i56
	assign leaf[860] = !f[369] && f[402] && !f[526] && f[318]; // c3t563i56
	assign leaf[861] = !f[369] && f[402] && f[526] && !f[126]; // c3t563i56
	assign leaf[862] = !f[369] && f[402] && f[526] && f[126]; // c3t563i56
	assign leaf[863] = f[369] && !f[544] && !f[217] && !f[293]; // c3t563i56
	assign leaf[864] = f[369] && !f[544] && !f[217] && f[293]; // c3t563i56
	assign leaf[865] = f[369] && !f[544] && f[217]; // c3t563i56
	assign leaf[866] = f[369] && f[544] && !f[234]; // c3t563i56
	assign leaf[867] = f[369] && f[544] && f[234]; // c3t563i56
	assign leaf[868] = !f[708] && !f[357] && !f[190] && !f[649]; // c3t573i57
	assign leaf[869] = !f[708] && !f[357] && !f[190] && f[649]; // c3t573i57
	assign leaf[870] = !f[708] && !f[357] && f[190] && !f[355]; // c3t573i57
	assign leaf[871] = !f[708] && !f[357] && f[190] && f[355]; // c3t573i57
	assign leaf[872] = !f[708] && f[357] && !f[266] && !f[160]; // c3t573i57
	assign leaf[873] = !f[708] && f[357] && !f[266] && f[160]; // c3t573i57
	assign leaf[874] = !f[708] && f[357] && f[266] && !f[187]; // c3t573i57
	assign leaf[875] = !f[708] && f[357] && f[266] && f[187]; // c3t573i57
	assign leaf[876] = f[708] && !f[599] && !f[518] && !f[244]; // c3t573i57
	assign leaf[877] = f[708] && !f[599] && !f[518] && f[244]; // c3t573i57
	assign leaf[878] = f[708] && !f[599] && f[518]; // c3t573i57
	assign leaf[879] = f[708] && f[599] && !f[602]; // c3t573i57
	assign leaf[880] = f[708] && f[599] && f[602]; // c3t573i57
	assign leaf[881] = !f[384] && !f[495] && !f[293] && !f[298]; // c3t583i58
	assign leaf[882] = !f[384] && !f[495] && !f[293] && f[298]; // c3t583i58
	assign leaf[883] = !f[384] && !f[495] && f[293] && !f[319]; // c3t583i58
	assign leaf[884] = !f[384] && !f[495] && f[293] && f[319]; // c3t583i58
	assign leaf[885] = !f[384] && f[495] && !f[442] && !f[435]; // c3t583i58
	assign leaf[886] = !f[384] && f[495] && !f[442] && f[435]; // c3t583i58
	assign leaf[887] = !f[384] && f[495] && f[442]; // c3t583i58
	assign leaf[888] = f[384] && !f[438] && !f[353] && !f[537]; // c3t583i58
	assign leaf[889] = f[384] && !f[438] && !f[353] && f[537]; // c3t583i58
	assign leaf[890] = f[384] && !f[438] && f[353] && !f[211]; // c3t583i58
	assign leaf[891] = f[384] && !f[438] && f[353] && f[211]; // c3t583i58
	assign leaf[892] = f[384] && f[438] && !f[517] && !f[327]; // c3t583i58
	assign leaf[893] = f[384] && f[438] && !f[517] && f[327]; // c3t583i58
	assign leaf[894] = f[384] && f[438] && f[517] && !f[126]; // c3t583i58
	assign leaf[895] = f[384] && f[438] && f[517] && f[126]; // c3t583i58
	assign leaf[896] = !f[492] && !f[547] && !f[517] && !f[407]; // c3t593i59
	assign leaf[897] = !f[492] && !f[547] && !f[517] && f[407]; // c3t593i59
	assign leaf[898] = !f[492] && !f[547] && f[517] && !f[572]; // c3t593i59
	assign leaf[899] = !f[492] && !f[547] && f[517] && f[572]; // c3t593i59
	assign leaf[900] = !f[492] && f[547] && !f[409] && !f[581]; // c3t593i59
	assign leaf[901] = !f[492] && f[547] && !f[409] && f[581]; // c3t593i59
	assign leaf[902] = !f[492] && f[547] && f[409] && !f[516]; // c3t593i59
	assign leaf[903] = !f[492] && f[547] && f[409] && f[516]; // c3t593i59
	assign leaf[904] = f[492] && !f[438] && !f[493] && !f[293]; // c3t593i59
	assign leaf[905] = f[492] && !f[438] && !f[493] && f[293]; // c3t593i59
	assign leaf[906] = f[492] && !f[438] && f[493] && !f[355]; // c3t593i59
	assign leaf[907] = f[492] && !f[438] && f[493] && f[355]; // c3t593i59
	assign leaf[908] = f[492] && f[438] && !f[295] && !f[564]; // c3t593i59
	assign leaf[909] = f[492] && f[438] && !f[295] && f[564]; // c3t593i59
	assign leaf[910] = f[492] && f[438] && f[295] && !f[155]; // c3t593i59
	assign leaf[911] = f[492] && f[438] && f[295] && f[155]; // c3t593i59
	assign leaf[912] = !f[429] && !f[127] && !f[209] && !f[173]; // c3t603i60
	assign leaf[913] = !f[429] && !f[127] && !f[209] && f[173]; // c3t603i60
	assign leaf[914] = !f[429] && !f[127] && f[209] && !f[320]; // c3t603i60
	assign leaf[915] = !f[429] && !f[127] && f[209] && f[320]; // c3t603i60
	assign leaf[916] = !f[429] && f[127] && !f[459] && !f[235]; // c3t603i60
	assign leaf[917] = !f[429] && f[127] && !f[459] && f[235]; // c3t603i60
	assign leaf[918] = !f[429] && f[127] && f[459] && !f[652]; // c3t603i60
	assign leaf[919] = !f[429] && f[127] && f[459] && f[652]; // c3t603i60
	assign leaf[920] = f[429] && !f[544] && !f[513] && !f[553]; // c3t603i60
	assign leaf[921] = f[429] && !f[544] && !f[513] && f[553]; // c3t603i60
	assign leaf[922] = f[429] && !f[544] && f[513] && !f[130]; // c3t603i60
	assign leaf[923] = f[429] && !f[544] && f[513] && f[130]; // c3t603i60
	assign leaf[924] = f[429] && f[544] && !f[687] && !f[549]; // c3t603i60
	assign leaf[925] = f[429] && f[544] && !f[687] && f[549]; // c3t603i60
	assign leaf[926] = f[429] && f[544] && f[687] && !f[327]; // c3t603i60
	assign leaf[927] = f[429] && f[544] && f[687] && f[327]; // c3t603i60
	assign leaf[928] = !f[384] && !f[358] && !f[328] && !f[190]; // c3t613i61
	assign leaf[929] = !f[384] && !f[358] && !f[328] && f[190]; // c3t613i61
	assign leaf[930] = !f[384] && !f[358] && f[328] && !f[241]; // c3t613i61
	assign leaf[931] = !f[384] && !f[358] && f[328] && f[241]; // c3t613i61
	assign leaf[932] = !f[384] && f[358]; // c3t613i61
	assign leaf[933] = f[384] && !f[266] && !f[131] && !f[461]; // c3t613i61
	assign leaf[934] = f[384] && !f[266] && !f[131] && f[461]; // c3t613i61
	assign leaf[935] = f[384] && !f[266] && f[131] && !f[236]; // c3t613i61
	assign leaf[936] = f[384] && !f[266] && f[131] && f[236]; // c3t613i61
	assign leaf[937] = f[384] && f[266] && !f[122] && !f[298]; // c3t613i61
	assign leaf[938] = f[384] && f[266] && !f[122] && f[298]; // c3t613i61
	assign leaf[939] = f[384] && f[266] && f[122] && !f[261]; // c3t613i61
	assign leaf[940] = f[384] && f[266] && f[122] && f[261]; // c3t613i61
	assign leaf[941] = !f[705] && !f[386] && !f[346] && !f[372]; // c3t623i62
	assign leaf[942] = !f[705] && !f[386] && !f[346] && f[372]; // c3t623i62
	assign leaf[943] = !f[705] && !f[386] && f[346] && !f[321]; // c3t623i62
	assign leaf[944] = !f[705] && !f[386] && f[346] && f[321]; // c3t623i62
	assign leaf[945] = !f[705] && f[386] && !f[152] && !f[508]; // c3t623i62
	assign leaf[946] = !f[705] && f[386] && !f[152] && f[508]; // c3t623i62
	assign leaf[947] = !f[705] && f[386] && f[152] && !f[237]; // c3t623i62
	assign leaf[948] = !f[705] && f[386] && f[152] && f[237]; // c3t623i62
	assign leaf[949] = f[705]; // c3t623i62
	assign leaf[950] = !f[707] && !f[571] && !f[546] && !f[490]; // c3t633i63
	assign leaf[951] = !f[707] && !f[571] && !f[546] && f[490]; // c3t633i63
	assign leaf[952] = !f[707] && !f[571] && f[546] && !f[492]; // c3t633i63
	assign leaf[953] = !f[707] && !f[571] && f[546] && f[492]; // c3t633i63
	assign leaf[954] = !f[707] && f[571] && !f[596] && !f[580]; // c3t633i63
	assign leaf[955] = !f[707] && f[571] && !f[596] && f[580]; // c3t633i63
	assign leaf[956] = !f[707] && f[571] && f[596] && !f[519]; // c3t633i63
	assign leaf[957] = !f[707] && f[571] && f[596] && f[519]; // c3t633i63
	assign leaf[958] = f[707] && !f[267]; // c3t633i63
	assign leaf[959] = f[707] && f[267] && !f[571]; // c3t633i63
	assign leaf[960] = f[707] && f[267] && f[571]; // c3t633i63
	assign leaf[961] = !f[346] && !f[290] && !f[292] && !f[376]; // c3t643i64
	assign leaf[962] = !f[346] && !f[290] && !f[292] && f[376]; // c3t643i64
	assign leaf[963] = !f[346] && !f[290] && f[292] && !f[266]; // c3t643i64
	assign leaf[964] = !f[346] && !f[290] && f[292] && f[266]; // c3t643i64
	assign leaf[965] = !f[346] && f[290] && !f[320] && !f[129]; // c3t643i64
	assign leaf[966] = !f[346] && f[290] && !f[320] && f[129]; // c3t643i64
	assign leaf[967] = !f[346] && f[290] && f[320] && !f[238]; // c3t643i64
	assign leaf[968] = !f[346] && f[290] && f[320] && f[238]; // c3t643i64
	assign leaf[969] = f[346] && !f[321] && !f[403] && !f[327]; // c3t643i64
	assign leaf[970] = f[346] && !f[321] && !f[403] && f[327]; // c3t643i64
	assign leaf[971] = f[346] && !f[321] && f[403] && !f[636]; // c3t643i64
	assign leaf[972] = f[346] && !f[321] && f[403] && f[636]; // c3t643i64
	assign leaf[973] = f[346] && f[321] && !f[289] && !f[152]; // c3t643i64
	assign leaf[974] = f[346] && f[321] && !f[289] && f[152]; // c3t643i64
	assign leaf[975] = f[346] && f[321] && f[289] && !f[627]; // c3t643i64
	assign leaf[976] = f[346] && f[321] && f[289] && f[627]; // c3t643i64
	assign leaf[977] = !f[399] && !f[740] && !f[626] && !f[600]; // c3t653i65
	assign leaf[978] = !f[399] && !f[740] && !f[626] && f[600]; // c3t653i65
	assign leaf[979] = !f[399] && !f[740] && f[626] && !f[629]; // c3t653i65
	assign leaf[980] = !f[399] && !f[740] && f[626] && f[629]; // c3t653i65
	assign leaf[981] = !f[399] && f[740]; // c3t653i65
	assign leaf[982] = f[399] && !f[411] && !f[186] && !f[454]; // c3t653i65
	assign leaf[983] = f[399] && !f[411] && !f[186] && f[454]; // c3t653i65
	assign leaf[984] = f[399] && !f[411] && f[186] && !f[682]; // c3t653i65
	assign leaf[985] = f[399] && !f[411] && f[186] && f[682]; // c3t653i65
	assign leaf[986] = f[399] && f[411] && !f[294] && !f[408]; // c3t653i65
	assign leaf[987] = f[399] && f[411] && !f[294] && f[408]; // c3t653i65
	assign leaf[988] = f[399] && f[411] && f[294] && !f[317]; // c3t653i65
	assign leaf[989] = f[399] && f[411] && f[294] && f[317]; // c3t653i65
	assign leaf[990] = !f[429] && !f[213] && !f[713] && !f[458]; // c3t663i66
	assign leaf[991] = !f[429] && !f[213] && !f[713] && f[458]; // c3t663i66
	assign leaf[992] = !f[429] && !f[213] && f[713] && !f[323]; // c3t663i66
	assign leaf[993] = !f[429] && !f[213] && f[713] && f[323]; // c3t663i66
	assign leaf[994] = !f[429] && f[213] && !f[126] && !f[570]; // c3t663i66
	assign leaf[995] = !f[429] && f[213] && !f[126] && f[570]; // c3t663i66
	assign leaf[996] = !f[429] && f[213] && f[126] && !f[487]; // c3t663i66
	assign leaf[997] = !f[429] && f[213] && f[126] && f[487]; // c3t663i66
	assign leaf[998] = f[429] && !f[459] && !f[483] && !f[485]; // c3t663i66
	assign leaf[999] = f[429] && !f[459] && !f[483] && f[485]; // c3t663i66
	assign leaf[1000] = f[429] && !f[459] && f[483] && !f[498]; // c3t663i66
	assign leaf[1001] = f[429] && !f[459] && f[483] && f[498]; // c3t663i66
	assign leaf[1002] = f[429] && f[459] && !f[346] && !f[580]; // c3t663i66
	assign leaf[1003] = f[429] && f[459] && !f[346] && f[580]; // c3t663i66
	assign leaf[1004] = f[429] && f[459] && f[346] && !f[182]; // c3t663i66
	assign leaf[1005] = f[429] && f[459] && f[346] && f[182]; // c3t663i66
	assign leaf[1006] = !f[386] && !f[537] && !f[570] && !f[460]; // c3t673i67
	assign leaf[1007] = !f[386] && !f[537] && !f[570] && f[460]; // c3t673i67
	assign leaf[1008] = !f[386] && !f[537] && f[570] && !f[600]; // c3t673i67
	assign leaf[1009] = !f[386] && !f[537] && f[570] && f[600]; // c3t673i67
	assign leaf[1010] = !f[386] && f[537] && !f[302] && !f[602]; // c3t673i67
	assign leaf[1011] = !f[386] && f[537] && !f[302] && f[602]; // c3t673i67
	assign leaf[1012] = !f[386] && f[537] && f[302] && !f[483]; // c3t673i67
	assign leaf[1013] = !f[386] && f[537] && f[302] && f[483]; // c3t673i67
	assign leaf[1014] = f[386] && !f[355]; // c3t673i67
	assign leaf[1015] = f[386] && f[355] && !f[580] && !f[185]; // c3t673i67
	assign leaf[1016] = f[386] && f[355] && !f[580] && f[185]; // c3t673i67
	assign leaf[1017] = f[386] && f[355] && f[580] && !f[259]; // c3t673i67
	assign leaf[1018] = f[386] && f[355] && f[580] && f[259]; // c3t673i67
	assign leaf[1019] = !f[682] && !f[626] && !f[602] && !f[714]; // c3t683i68
	assign leaf[1020] = !f[682] && !f[626] && !f[602] && f[714]; // c3t683i68
	assign leaf[1021] = !f[682] && !f[626] && f[602] && !f[598]; // c3t683i68
	assign leaf[1022] = !f[682] && !f[626] && f[602] && f[598]; // c3t683i68
	assign leaf[1023] = !f[682] && f[626] && !f[431] && !f[207]; // c3t683i68
	assign leaf[1024] = !f[682] && f[626] && !f[431] && f[207]; // c3t683i68
	assign leaf[1025] = !f[682] && f[626] && f[431] && !f[485]; // c3t683i68
	assign leaf[1026] = !f[682] && f[626] && f[431] && f[485]; // c3t683i68
	assign leaf[1027] = f[682] && !f[541] && !f[320] && !f[602]; // c3t683i68
	assign leaf[1028] = f[682] && !f[541] && !f[320] && f[602]; // c3t683i68
	assign leaf[1029] = f[682] && !f[541] && f[320] && !f[598]; // c3t683i68
	assign leaf[1030] = f[682] && !f[541] && f[320] && f[598]; // c3t683i68
	assign leaf[1031] = f[682] && f[541] && !f[514] && !f[299]; // c3t683i68
	assign leaf[1032] = f[682] && f[541] && !f[514] && f[299]; // c3t683i68
	assign leaf[1033] = f[682] && f[541] && f[514] && !f[407]; // c3t683i68
	assign leaf[1034] = f[682] && f[541] && f[514] && f[407]; // c3t683i68
	assign leaf[1035] = !f[434] && !f[321] && !f[96] && !f[351]; // c3t693i69
	assign leaf[1036] = !f[434] && !f[321] && !f[96] && f[351]; // c3t693i69
	assign leaf[1037] = !f[434] && !f[321] && f[96] && !f[549]; // c3t693i69
	assign leaf[1038] = !f[434] && !f[321] && f[96] && f[549]; // c3t693i69
	assign leaf[1039] = !f[434] && f[321] && !f[347] && !f[436]; // c3t693i69
	assign leaf[1040] = !f[434] && f[321] && !f[347] && f[436]; // c3t693i69
	assign leaf[1041] = !f[434] && f[321] && f[347] && !f[288]; // c3t693i69
	assign leaf[1042] = !f[434] && f[321] && f[347] && f[288]; // c3t693i69
	assign leaf[1043] = f[434] && !f[208] && !f[461] && !f[406]; // c3t693i69
	assign leaf[1044] = f[434] && !f[208] && !f[461] && f[406]; // c3t693i69
	assign leaf[1045] = f[434] && !f[208] && f[461] && !f[606]; // c3t693i69
	assign leaf[1046] = f[434] && !f[208] && f[461] && f[606]; // c3t693i69
	assign leaf[1047] = f[434] && f[208] && !f[572] && !f[516]; // c3t693i69
	assign leaf[1048] = f[434] && f[208] && !f[572] && f[516]; // c3t693i69
	assign leaf[1049] = f[434] && f[208] && f[572] && !f[489]; // c3t693i69
	assign leaf[1050] = f[434] && f[208] && f[572] && f[489]; // c3t693i69
	assign leaf[1051] = !f[402] && !f[709] && !f[266] && !f[378]; // c3t703i70
	assign leaf[1052] = !f[402] && !f[709] && !f[266] && f[378]; // c3t703i70
	assign leaf[1053] = !f[402] && !f[709] && f[266] && !f[160]; // c3t703i70
	assign leaf[1054] = !f[402] && !f[709] && f[266] && f[160]; // c3t703i70
	assign leaf[1055] = !f[402] && f[709] && !f[320] && !f[630]; // c3t703i70
	assign leaf[1056] = !f[402] && f[709] && !f[320] && f[630]; // c3t703i70
	assign leaf[1057] = !f[402] && f[709] && f[320]; // c3t703i70
	assign leaf[1058] = f[402] && !f[512] && !f[482] && !f[349]; // c3t703i70
	assign leaf[1059] = f[402] && !f[512] && !f[482] && f[349]; // c3t703i70
	assign leaf[1060] = f[402] && !f[512] && f[482] && !f[434]; // c3t703i70
	assign leaf[1061] = f[402] && !f[512] && f[482] && f[434]; // c3t703i70
	assign leaf[1062] = f[402] && f[512] && !f[457] && !f[269]; // c3t703i70
	assign leaf[1063] = f[402] && f[512] && !f[457] && f[269]; // c3t703i70
	assign leaf[1064] = f[402] && f[512] && f[457] && !f[454]; // c3t703i70
	assign leaf[1065] = f[402] && f[512] && f[457] && f[454]; // c3t703i70
	assign leaf[1066] = !f[712] && !f[718] && !f[626] && !f[683]; // c3t713i71
	assign leaf[1067] = !f[712] && !f[718] && !f[626] && f[683]; // c3t713i71
	assign leaf[1068] = !f[712] && !f[718] && f[626] && !f[426]; // c3t713i71
	assign leaf[1069] = !f[712] && !f[718] && f[626] && f[426]; // c3t713i71
	assign leaf[1070] = !f[712] && f[718] && !f[489] && !f[459]; // c3t713i71
	assign leaf[1071] = !f[712] && f[718] && !f[489] && f[459]; // c3t713i71
	assign leaf[1072] = !f[712] && f[718] && f[489] && !f[493]; // c3t713i71
	assign leaf[1073] = !f[712] && f[718] && f[489] && f[493]; // c3t713i71
	assign leaf[1074] = f[712] && !f[375] && !f[409] && !f[433]; // c3t713i71
	assign leaf[1075] = f[712] && !f[375] && !f[409] && f[433]; // c3t713i71
	assign leaf[1076] = f[712] && !f[375] && f[409] && !f[430]; // c3t713i71
	assign leaf[1077] = f[712] && !f[375] && f[409] && f[430]; // c3t713i71
	assign leaf[1078] = f[712] && f[375] && !f[322] && !f[263]; // c3t713i71
	assign leaf[1079] = f[712] && f[375] && !f[322] && f[263]; // c3t713i71
	assign leaf[1080] = f[712] && f[375] && f[322] && !f[319]; // c3t713i71
	assign leaf[1081] = f[712] && f[375] && f[322] && f[319]; // c3t713i71
	assign leaf[1082] = !f[373] && !f[689] && !f[740] && !f[715]; // c3t723i72
	assign leaf[1083] = !f[373] && !f[689] && !f[740] && f[715]; // c3t723i72
	assign leaf[1084] = !f[373] && !f[689] && f[740]; // c3t723i72
	assign leaf[1085] = !f[373] && f[689] && !f[575] && !f[519]; // c3t723i72
	assign leaf[1086] = !f[373] && f[689] && !f[575] && f[519]; // c3t723i72
	assign leaf[1087] = !f[373] && f[689] && f[575] && !f[492]; // c3t723i72
	assign leaf[1088] = !f[373] && f[689] && f[575] && f[492]; // c3t723i72
	assign leaf[1089] = f[373] && !f[320] && !f[264] && !f[233]; // c3t723i72
	assign leaf[1090] = f[373] && !f[320] && !f[264] && f[233]; // c3t723i72
	assign leaf[1091] = f[373] && !f[320] && f[264] && !f[239]; // c3t723i72
	assign leaf[1092] = f[373] && !f[320] && f[264] && f[239]; // c3t723i72
	assign leaf[1093] = f[373] && f[320] && !f[298] && !f[216]; // c3t723i72
	assign leaf[1094] = f[373] && f[320] && !f[298] && f[216]; // c3t723i72
	assign leaf[1095] = f[373] && f[320] && f[298] && !f[155]; // c3t723i72
	assign leaf[1096] = f[373] && f[320] && f[298] && f[155]; // c3t723i72
	assign leaf[1097] = !f[331] && !f[676] && !f[479] && !f[604]; // c3t733i73
	assign leaf[1098] = !f[331] && !f[676] && !f[479] && f[604]; // c3t733i73
	assign leaf[1099] = !f[331] && !f[676] && f[479] && !f[426]; // c3t733i73
	assign leaf[1100] = !f[331] && !f[676] && f[479] && f[426]; // c3t733i73
	assign leaf[1101] = !f[331] && f[676]; // c3t733i73
	assign leaf[1102] = f[331] && !f[234]; // c3t733i73
	assign leaf[1103] = f[331] && f[234]; // c3t733i73
	assign leaf[1104] = !f[120] && !f[269] && !f[296] && !f[513]; // c3t743i74
	assign leaf[1105] = !f[120] && !f[269] && !f[296] && f[513]; // c3t743i74
	assign leaf[1106] = !f[120] && !f[269] && f[296] && !f[129]; // c3t743i74
	assign leaf[1107] = !f[120] && !f[269] && f[296] && f[129]; // c3t743i74
	assign leaf[1108] = !f[120] && f[269] && !f[101] && !f[378]; // c3t743i74
	assign leaf[1109] = !f[120] && f[269] && !f[101] && f[378]; // c3t743i74
	assign leaf[1110] = !f[120] && f[269] && f[101] && !f[579]; // c3t743i74
	assign leaf[1111] = !f[120] && f[269] && f[101] && f[579]; // c3t743i74
	assign leaf[1112] = f[120] && !f[630]; // c3t743i74
	assign leaf[1113] = f[120] && f[630] && !f[458] && !f[292]; // c3t743i74
	assign leaf[1114] = f[120] && f[630] && !f[458] && f[292]; // c3t743i74
	assign leaf[1115] = f[120] && f[630] && f[458]; // c3t743i74
	assign leaf[1116] = !f[712] && !f[313] && !f[202] && !f[258]; // c3t753i75
	assign leaf[1117] = !f[712] && !f[313] && !f[202] && f[258]; // c3t753i75
	assign leaf[1118] = !f[712] && !f[313] && f[202] && !f[576]; // c3t753i75
	assign leaf[1119] = !f[712] && !f[313] && f[202] && f[576]; // c3t753i75
	assign leaf[1120] = !f[712] && f[313] && !f[525] && !f[685]; // c3t753i75
	assign leaf[1121] = !f[712] && f[313] && !f[525] && f[685]; // c3t753i75
	assign leaf[1122] = !f[712] && f[313] && f[525] && !f[397]; // c3t753i75
	assign leaf[1123] = !f[712] && f[313] && f[525] && f[397]; // c3t753i75
	assign leaf[1124] = f[712] && !f[684] && !f[178]; // c3t753i75
	assign leaf[1125] = f[712] && !f[684] && f[178]; // c3t753i75
	assign leaf[1126] = f[712] && f[684] && !f[576] && !f[356]; // c3t753i75
	assign leaf[1127] = f[712] && f[684] && !f[576] && f[356]; // c3t753i75
	assign leaf[1128] = f[712] && f[684] && f[576] && !f[299]; // c3t753i75
	assign leaf[1129] = f[712] && f[684] && f[576] && f[299]; // c3t753i75
	assign leaf[1130] = !f[708] && !f[466] && !f[718] && !f[200]; // c3t763i76
	assign leaf[1131] = !f[708] && !f[466] && !f[718] && f[200]; // c3t763i76
	assign leaf[1132] = !f[708] && !f[466] && f[718] && !f[213]; // c3t763i76
	assign leaf[1133] = !f[708] && !f[466] && f[718] && f[213]; // c3t763i76
	assign leaf[1134] = !f[708] && f[466] && !f[355] && !f[403]; // c3t763i76
	assign leaf[1135] = !f[708] && f[466] && !f[355] && f[403]; // c3t763i76
	assign leaf[1136] = !f[708] && f[466] && f[355] && !f[543]; // c3t763i76
	assign leaf[1137] = !f[708] && f[466] && f[355] && f[543]; // c3t763i76
	assign leaf[1138] = f[708] && !f[599] && !f[491]; // c3t763i76
	assign leaf[1139] = f[708] && !f[599] && f[491]; // c3t763i76
	assign leaf[1140] = f[708] && f[599]; // c3t763i76
	assign leaf[1141] = !f[427] && !f[651] && !f[712] && !f[626]; // c3t773i77
	assign leaf[1142] = !f[427] && !f[651] && !f[712] && f[626]; // c3t773i77
	assign leaf[1143] = !f[427] && !f[651] && f[712] && !f[488]; // c3t773i77
	assign leaf[1144] = !f[427] && !f[651] && f[712] && f[488]; // c3t773i77
	assign leaf[1145] = !f[427] && f[651] && !f[542] && !f[461]; // c3t773i77
	assign leaf[1146] = !f[427] && f[651] && !f[542] && f[461]; // c3t773i77
	assign leaf[1147] = !f[427] && f[651] && f[542] && !f[656]; // c3t773i77
	assign leaf[1148] = !f[427] && f[651] && f[542] && f[656]; // c3t773i77
	assign leaf[1149] = f[427] && !f[436] && !f[236] && !f[295]; // c3t773i77
	assign leaf[1150] = f[427] && !f[436] && !f[236] && f[295]; // c3t773i77
	assign leaf[1151] = f[427] && !f[436] && f[236] && !f[597]; // c3t773i77
	assign leaf[1152] = f[427] && !f[436] && f[236] && f[597]; // c3t773i77
	assign leaf[1153] = f[427] && f[436] && !f[580] && !f[568]; // c3t773i77
	assign leaf[1154] = f[427] && f[436] && !f[580] && f[568]; // c3t773i77
	assign leaf[1155] = f[427] && f[436] && f[580] && !f[658]; // c3t773i77
	assign leaf[1156] = f[427] && f[436] && f[580] && f[658]; // c3t773i77
	assign leaf[1157] = !f[384] && !f[487] && !f[124] && !f[554]; // c3t783i78
	assign leaf[1158] = !f[384] && !f[487] && !f[124] && f[554]; // c3t783i78
	assign leaf[1159] = !f[384] && !f[487] && f[124] && !f[207]; // c3t783i78
	assign leaf[1160] = !f[384] && !f[487] && f[124] && f[207]; // c3t783i78
	assign leaf[1161] = !f[384] && f[487] && !f[570] && !f[294]; // c3t783i78
	assign leaf[1162] = !f[384] && f[487] && !f[570] && f[294]; // c3t783i78
	assign leaf[1163] = !f[384] && f[487] && f[570] && !f[460]; // c3t783i78
	assign leaf[1164] = !f[384] && f[487] && f[570] && f[460]; // c3t783i78
	assign leaf[1165] = f[384] && !f[295] && !f[439] && !f[496]; // c3t783i78
	assign leaf[1166] = f[384] && !f[295] && !f[439] && f[496]; // c3t783i78
	assign leaf[1167] = f[384] && !f[295] && f[439] && !f[158]; // c3t783i78
	assign leaf[1168] = f[384] && !f[295] && f[439] && f[158]; // c3t783i78
	assign leaf[1169] = f[384] && f[295] && !f[239] && !f[261]; // c3t783i78
	assign leaf[1170] = f[384] && f[295] && !f[239] && f[261]; // c3t783i78
	assign leaf[1171] = f[384] && f[295] && f[239] && !f[126]; // c3t783i78
	assign leaf[1172] = f[384] && f[295] && f[239] && f[126]; // c3t783i78
	assign leaf[1173] = !f[346] && !f[433] && !f[462] && !f[314]; // c3t793i79
	assign leaf[1174] = !f[346] && !f[433] && !f[462] && f[314]; // c3t793i79
	assign leaf[1175] = !f[346] && !f[433] && f[462] && !f[298]; // c3t793i79
	assign leaf[1176] = !f[346] && !f[433] && f[462] && f[298]; // c3t793i79
	assign leaf[1177] = !f[346] && f[433] && !f[321] && !f[372]; // c3t793i79
	assign leaf[1178] = !f[346] && f[433] && !f[321] && f[372]; // c3t793i79
	assign leaf[1179] = !f[346] && f[433] && f[321] && !f[180]; // c3t793i79
	assign leaf[1180] = !f[346] && f[433] && f[321] && f[180]; // c3t793i79
	assign leaf[1181] = f[346] && !f[470] && !f[375] && !f[378]; // c3t793i79
	assign leaf[1182] = f[346] && !f[470] && !f[375] && f[378]; // c3t793i79
	assign leaf[1183] = f[346] && !f[470] && f[375] && !f[289]; // c3t793i79
	assign leaf[1184] = f[346] && !f[470] && f[375] && f[289]; // c3t793i79
	assign leaf[1185] = f[346] && f[470] && !f[463] && !f[410]; // c3t793i79
	assign leaf[1186] = f[346] && f[470] && !f[463] && f[410]; // c3t793i79
	assign leaf[1187] = f[346] && f[470] && f[463]; // c3t793i79
	assign leaf[1188] = !f[209] && !f[265] && !f[261] && !f[235]; // c3t803i80
	assign leaf[1189] = !f[209] && !f[265] && !f[261] && f[235]; // c3t803i80
	assign leaf[1190] = !f[209] && !f[265] && f[261] && !f[470]; // c3t803i80
	assign leaf[1191] = !f[209] && !f[265] && f[261] && f[470]; // c3t803i80
	assign leaf[1192] = !f[209] && f[265] && !f[126] && !f[321]; // c3t803i80
	assign leaf[1193] = !f[209] && f[265] && !f[126] && f[321]; // c3t803i80
	assign leaf[1194] = !f[209] && f[265] && f[126] && !f[239]; // c3t803i80
	assign leaf[1195] = !f[209] && f[265] && f[126] && f[239]; // c3t803i80
	assign leaf[1196] = f[209] && !f[98] && !f[435] && !f[315]; // c3t803i80
	assign leaf[1197] = f[209] && !f[98] && !f[435] && f[315]; // c3t803i80
	assign leaf[1198] = f[209] && !f[98] && f[435] && !f[379]; // c3t803i80
	assign leaf[1199] = f[209] && !f[98] && f[435] && f[379]; // c3t803i80
	assign leaf[1200] = f[209] && f[98] && !f[123]; // c3t803i80
	assign leaf[1201] = f[209] && f[98] && f[123]; // c3t803i80
	assign leaf[1202] = !f[429] && !f[96] && !f[178] && !f[241]; // c3t813i81
	assign leaf[1203] = !f[429] && !f[96] && !f[178] && f[241]; // c3t813i81
	assign leaf[1204] = !f[429] && !f[96] && f[178] && !f[261]; // c3t813i81
	assign leaf[1205] = !f[429] && !f[96] && f[178] && f[261]; // c3t813i81
	assign leaf[1206] = !f[429] && f[96] && !f[266] && !f[579]; // c3t813i81
	assign leaf[1207] = !f[429] && f[96] && !f[266] && f[579]; // c3t813i81
	assign leaf[1208] = !f[429] && f[96] && f[266] && !f[151]; // c3t813i81
	assign leaf[1209] = !f[429] && f[96] && f[266] && f[151]; // c3t813i81
	assign leaf[1210] = f[429] && !f[511] && !f[376] && !f[437]; // c3t813i81
	assign leaf[1211] = f[429] && !f[511] && !f[376] && f[437]; // c3t813i81
	assign leaf[1212] = f[429] && !f[511] && f[376] && !f[513]; // c3t813i81
	assign leaf[1213] = f[429] && !f[511] && f[376] && f[513]; // c3t813i81
	assign leaf[1214] = f[429] && f[511] && !f[542] && !f[434]; // c3t813i81
	assign leaf[1215] = f[429] && f[511] && !f[542] && f[434]; // c3t813i81
	assign leaf[1216] = f[429] && f[511] && f[542] && !f[181]; // c3t813i81
	assign leaf[1217] = f[429] && f[511] && f[542] && f[181]; // c3t813i81
	assign leaf[1218] = !f[705] && !f[358] && !f[330] && !f[357]; // c3t823i82
	assign leaf[1219] = !f[705] && !f[358] && !f[330] && f[357]; // c3t823i82
	assign leaf[1220] = !f[705] && !f[358] && f[330] && !f[321]; // c3t823i82
	assign leaf[1221] = !f[705] && !f[358] && f[330] && f[321]; // c3t823i82
	assign leaf[1222] = !f[705] && f[358] && !f[595]; // c3t823i82
	assign leaf[1223] = !f[705] && f[358] && f[595] && !f[576]; // c3t823i82
	assign leaf[1224] = !f[705] && f[358] && f[595] && f[576]; // c3t823i82
	assign leaf[1225] = f[705]; // c3t823i82
	assign leaf[1226] = !f[377] && !f[324] && !f[436] && !f[321]; // c3t833i83
	assign leaf[1227] = !f[377] && !f[324] && !f[436] && f[321]; // c3t833i83
	assign leaf[1228] = !f[377] && !f[324] && f[436] && !f[539]; // c3t833i83
	assign leaf[1229] = !f[377] && !f[324] && f[436] && f[539]; // c3t833i83
	assign leaf[1230] = !f[377] && f[324] && !f[436] && !f[547]; // c3t833i83
	assign leaf[1231] = !f[377] && f[324] && !f[436] && f[547]; // c3t833i83
	assign leaf[1232] = !f[377] && f[324] && f[436] && !f[604]; // c3t833i83
	assign leaf[1233] = !f[377] && f[324] && f[436] && f[604]; // c3t833i83
	assign leaf[1234] = f[377] && !f[181] && !f[126] && !f[263]; // c3t833i83
	assign leaf[1235] = f[377] && !f[181] && !f[126] && f[263]; // c3t833i83
	assign leaf[1236] = f[377] && !f[181] && f[126] && !f[436]; // c3t833i83
	assign leaf[1237] = f[377] && !f[181] && f[126] && f[436]; // c3t833i83
	assign leaf[1238] = f[377] && f[181] && !f[264] && !f[290]; // c3t833i83
	assign leaf[1239] = f[377] && f[181] && !f[264] && f[290]; // c3t833i83
	assign leaf[1240] = f[377] && f[181] && f[264] && !f[316]; // c3t833i83
	assign leaf[1241] = f[377] && f[181] && f[264] && f[316]; // c3t833i83
	assign leaf[1242] = !f[315] && !f[259] && !f[150] && !f[325]; // c3t843i84
	assign leaf[1243] = !f[315] && !f[259] && !f[150] && f[325]; // c3t843i84
	assign leaf[1244] = !f[315] && !f[259] && f[150] && !f[233]; // c3t843i84
	assign leaf[1245] = !f[315] && !f[259] && f[150] && f[233]; // c3t843i84
	assign leaf[1246] = !f[315] && f[259] && !f[375] && !f[572]; // c3t843i84
	assign leaf[1247] = !f[315] && f[259] && !f[375] && f[572]; // c3t843i84
	assign leaf[1248] = !f[315] && f[259] && f[375] && !f[149]; // c3t843i84
	assign leaf[1249] = !f[315] && f[259] && f[375] && f[149]; // c3t843i84
	assign leaf[1250] = f[315] && !f[345] && !f[399] && !f[433]; // c3t843i84
	assign leaf[1251] = f[315] && !f[345] && !f[399] && f[433]; // c3t843i84
	assign leaf[1252] = f[315] && !f[345] && f[399]; // c3t843i84
	assign leaf[1253] = f[315] && f[345] && !f[291] && !f[625]; // c3t843i84
	assign leaf[1254] = f[315] && f[345] && !f[291] && f[625]; // c3t843i84
	assign leaf[1255] = f[315] && f[345] && f[291] && !f[238]; // c3t843i84
	assign leaf[1256] = f[315] && f[345] && f[291] && f[238]; // c3t843i84
	assign leaf[1257] = !f[406] && !f[315] && !f[517] && !f[348]; // c3t853i85
	assign leaf[1258] = !f[406] && !f[315] && !f[517] && f[348]; // c3t853i85
	assign leaf[1259] = !f[406] && !f[315] && f[517] && !f[296]; // c3t853i85
	assign leaf[1260] = !f[406] && !f[315] && f[517] && f[296]; // c3t853i85
	assign leaf[1261] = !f[406] && f[315] && !f[438] && !f[327]; // c3t853i85
	assign leaf[1262] = !f[406] && f[315] && !f[438] && f[327]; // c3t853i85
	assign leaf[1263] = !f[406] && f[315] && f[438] && !f[489]; // c3t853i85
	assign leaf[1264] = !f[406] && f[315] && f[438] && f[489]; // c3t853i85
	assign leaf[1265] = f[406] && !f[604] && !f[608] && !f[547]; // c3t853i85
	assign leaf[1266] = f[406] && !f[604] && !f[608] && f[547]; // c3t853i85
	assign leaf[1267] = f[406] && !f[604] && f[608] && !f[235]; // c3t853i85
	assign leaf[1268] = f[406] && !f[604] && f[608] && f[235]; // c3t853i85
	assign leaf[1269] = f[406] && f[604] && !f[346] && !f[380]; // c3t853i85
	assign leaf[1270] = f[406] && f[604] && !f[346] && f[380]; // c3t853i85
	assign leaf[1271] = f[406] && f[604] && f[346] && !f[403]; // c3t853i85
	assign leaf[1272] = f[406] && f[604] && f[346] && f[403]; // c3t853i85
	assign leaf[1273] = !f[386] && !f[401] && !f[347] && !f[290]; // c3t863i86
	assign leaf[1274] = !f[386] && !f[401] && !f[347] && f[290]; // c3t863i86
	assign leaf[1275] = !f[386] && !f[401] && f[347] && !f[459]; // c3t863i86
	assign leaf[1276] = !f[386] && !f[401] && f[347] && f[459]; // c3t863i86
	assign leaf[1277] = !f[386] && f[401] && !f[509] && !f[442]; // c3t863i86
	assign leaf[1278] = !f[386] && f[401] && !f[509] && f[442]; // c3t863i86
	assign leaf[1279] = !f[386] && f[401] && f[509] && !f[454]; // c3t863i86
	assign leaf[1280] = !f[386] && f[401] && f[509] && f[454]; // c3t863i86
	assign leaf[1281] = f[386] && !f[499]; // c3t863i86
	assign leaf[1282] = f[386] && f[499] && !f[287]; // c3t863i86
	assign leaf[1283] = f[386] && f[499] && f[287]; // c3t863i86
	assign leaf[1284] = !f[707] && !f[344] && !f[270] && !f[187]; // c3t873i87
	assign leaf[1285] = !f[707] && !f[344] && !f[270] && f[187]; // c3t873i87
	assign leaf[1286] = !f[707] && !f[344] && f[270] && !f[293]; // c3t873i87
	assign leaf[1287] = !f[707] && !f[344] && f[270] && f[293]; // c3t873i87
	assign leaf[1288] = !f[707] && f[344] && !f[402] && !f[636]; // c3t873i87
	assign leaf[1289] = !f[707] && f[344] && !f[402] && f[636]; // c3t873i87
	assign leaf[1290] = !f[707] && f[344] && f[402] && !f[347]; // c3t873i87
	assign leaf[1291] = !f[707] && f[344] && f[402] && f[347]; // c3t873i87
	assign leaf[1292] = f[707] && !f[267]; // c3t873i87
	assign leaf[1293] = f[707] && f[267] && !f[493]; // c3t873i87
	assign leaf[1294] = f[707] && f[267] && f[493]; // c3t873i87
	assign leaf[1295] = !f[429] && !f[491] && !f[461] && !f[407]; // c3t883i88
	assign leaf[1296] = !f[429] && !f[491] && !f[461] && f[407]; // c3t883i88
	assign leaf[1297] = !f[429] && !f[491] && f[461] && !f[544]; // c3t883i88
	assign leaf[1298] = !f[429] && !f[491] && f[461] && f[544]; // c3t883i88
	assign leaf[1299] = !f[429] && f[491] && !f[461] && !f[233]; // c3t883i88
	assign leaf[1300] = !f[429] && f[491] && !f[461] && f[233]; // c3t883i88
	assign leaf[1301] = !f[429] && f[491] && f[461] && !f[662]; // c3t883i88
	assign leaf[1302] = !f[429] && f[491] && f[461] && f[662]; // c3t883i88
	assign leaf[1303] = f[429] && !f[526] && !f[544] && !f[266]; // c3t883i88
	assign leaf[1304] = f[429] && !f[526] && !f[544] && f[266]; // c3t883i88
	assign leaf[1305] = f[429] && !f[526] && f[544] && !f[267]; // c3t883i88
	assign leaf[1306] = f[429] && !f[526] && f[544] && f[267]; // c3t883i88
	assign leaf[1307] = f[429] && f[526] && !f[521] && !f[317]; // c3t883i88
	assign leaf[1308] = f[429] && f[526] && !f[521] && f[317]; // c3t883i88
	assign leaf[1309] = f[429] && f[526] && f[521]; // c3t883i88
	assign leaf[1310] = !f[549] && !f[487] && !f[458] && !f[346]; // c3t893i89
	assign leaf[1311] = !f[549] && !f[487] && !f[458] && f[346]; // c3t893i89
	assign leaf[1312] = !f[549] && !f[487] && f[458] && !f[209]; // c3t893i89
	assign leaf[1313] = !f[549] && !f[487] && f[458] && f[209]; // c3t893i89
	assign leaf[1314] = !f[549] && f[487] && !f[457] && !f[511]; // c3t893i89
	assign leaf[1315] = !f[549] && f[487] && !f[457] && f[511]; // c3t893i89
	assign leaf[1316] = !f[549] && f[487] && f[457] && !f[206]; // c3t893i89
	assign leaf[1317] = !f[549] && f[487] && f[457] && f[206]; // c3t893i89
	assign leaf[1318] = f[549] && !f[657] && !f[439] && !f[542]; // c3t893i89
	assign leaf[1319] = f[549] && !f[657] && !f[439] && f[542]; // c3t893i89
	assign leaf[1320] = f[549] && !f[657] && f[439] && !f[493]; // c3t893i89
	assign leaf[1321] = f[549] && !f[657] && f[439] && f[493]; // c3t893i89
	assign leaf[1322] = f[549] && f[657] && !f[384] && !f[687]; // c3t893i89
	assign leaf[1323] = f[549] && f[657] && !f[384] && f[687]; // c3t893i89
	assign leaf[1324] = f[549] && f[657] && f[384] && !f[522]; // c3t893i89
	assign leaf[1325] = f[549] && f[657] && f[384] && f[522]; // c3t893i89
	assign leaf[1326] = !f[492] && !f[547] && !f[517] && !f[322]; // c3t903i90
	assign leaf[1327] = !f[492] && !f[547] && !f[517] && f[322]; // c3t903i90
	assign leaf[1328] = !f[492] && !f[547] && f[517] && !f[572]; // c3t903i90
	assign leaf[1329] = !f[492] && !f[547] && f[517] && f[572]; // c3t903i90
	assign leaf[1330] = !f[492] && f[547] && !f[554] && !f[381]; // c3t903i90
	assign leaf[1331] = !f[492] && f[547] && !f[554] && f[381]; // c3t903i90
	assign leaf[1332] = !f[492] && f[547] && f[554] && !f[436]; // c3t903i90
	assign leaf[1333] = !f[492] && f[547] && f[554] && f[436]; // c3t903i90
	assign leaf[1334] = f[492] && !f[437] && !f[354] && !f[404]; // c3t903i90
	assign leaf[1335] = f[492] && !f[437] && !f[354] && f[404]; // c3t903i90
	assign leaf[1336] = f[492] && !f[437] && f[354] && !f[483]; // c3t903i90
	assign leaf[1337] = f[492] && !f[437] && f[354] && f[483]; // c3t903i90
	assign leaf[1338] = f[492] && f[437] && !f[625] && !f[274]; // c3t903i90
	assign leaf[1339] = f[492] && f[437] && !f[625] && f[274]; // c3t903i90
	assign leaf[1340] = f[492] && f[437] && f[625] && !f[154]; // c3t903i90
	assign leaf[1341] = f[492] && f[437] && f[625] && f[154]; // c3t903i90
	assign leaf[1342] = !f[427] && !f[705] && !f[591] && !f[218]; // c3t913i91
	assign leaf[1343] = !f[427] && !f[705] && !f[591] && f[218]; // c3t913i91
	assign leaf[1344] = !f[427] && !f[705] && f[591] && !f[159]; // c3t913i91
	assign leaf[1345] = !f[427] && !f[705] && f[591] && f[159]; // c3t913i91
	assign leaf[1346] = !f[427] && f[705]; // c3t913i91
	assign leaf[1347] = f[427] && !f[219] && !f[212] && !f[204]; // c3t913i91
	assign leaf[1348] = f[427] && !f[219] && !f[212] && f[204]; // c3t913i91
	assign leaf[1349] = f[427] && !f[219] && f[212] && !f[429]; // c3t913i91
	assign leaf[1350] = f[427] && !f[219] && f[212] && f[429]; // c3t913i91
	assign leaf[1351] = f[427] && f[219]; // c3t913i91
	assign leaf[1352] = !f[637] && !f[555] && !f[122] && !f[347]; // c3t923i92
	assign leaf[1353] = !f[637] && !f[555] && !f[122] && f[347]; // c3t923i92
	assign leaf[1354] = !f[637] && !f[555] && f[122] && !f[233]; // c3t923i92
	assign leaf[1355] = !f[637] && !f[555] && f[122] && f[233]; // c3t923i92
	assign leaf[1356] = !f[637] && f[555] && !f[320]; // c3t923i92
	assign leaf[1357] = !f[637] && f[555] && f[320] && !f[597]; // c3t923i92
	assign leaf[1358] = !f[637] && f[555] && f[320] && f[597]; // c3t923i92
	assign leaf[1359] = f[637] && !f[207] && !f[211]; // c3t923i92
	assign leaf[1360] = f[637] && !f[207] && f[211]; // c3t923i92
	assign leaf[1361] = f[637] && f[207] && !f[607] && !f[177]; // c3t923i92
	assign leaf[1362] = f[637] && f[207] && !f[607] && f[177]; // c3t923i92
	assign leaf[1363] = f[637] && f[207] && f[607] && !f[321]; // c3t923i92
	assign leaf[1364] = f[637] && f[207] && f[607] && f[321]; // c3t923i92
	assign leaf[1365] = !f[342] && !f[260] && !f[177] && !f[574]; // c3t933i93
	assign leaf[1366] = !f[342] && !f[260] && !f[177] && f[574]; // c3t933i93
	assign leaf[1367] = !f[342] && !f[260] && f[177] && !f[347]; // c3t933i93
	assign leaf[1368] = !f[342] && !f[260] && f[177] && f[347]; // c3t933i93
	assign leaf[1369] = !f[342] && f[260] && !f[289] && !f[347]; // c3t933i93
	assign leaf[1370] = !f[342] && f[260] && !f[289] && f[347]; // c3t933i93
	assign leaf[1371] = !f[342] && f[260] && f[289] && !f[236]; // c3t933i93
	assign leaf[1372] = !f[342] && f[260] && f[289] && f[236]; // c3t933i93
	assign leaf[1373] = f[342] && !f[323] && !f[355]; // c3t933i93
	assign leaf[1374] = f[342] && !f[323] && f[355] && !f[634]; // c3t933i93
	assign leaf[1375] = f[342] && !f[323] && f[355] && f[634]; // c3t933i93
	assign leaf[1376] = f[342] && f[323] && !f[525]; // c3t933i93
	assign leaf[1377] = f[342] && f[323] && f[525] && !f[270]; // c3t933i93
	assign leaf[1378] = f[342] && f[323] && f[525] && f[270]; // c3t933i93
	assign leaf[1379] = !f[406] && !f[517] && !f[325] && !f[217]; // c3t943i94
	assign leaf[1380] = !f[406] && !f[517] && !f[325] && f[217]; // c3t943i94
	assign leaf[1381] = !f[406] && !f[517] && f[325] && !f[437]; // c3t943i94
	assign leaf[1382] = !f[406] && !f[517] && f[325] && f[437]; // c3t943i94
	assign leaf[1383] = !f[406] && f[517] && !f[212] && !f[178]; // c3t943i94
	assign leaf[1384] = !f[406] && f[517] && !f[212] && f[178]; // c3t943i94
	assign leaf[1385] = !f[406] && f[517] && f[212] && !f[233]; // c3t943i94
	assign leaf[1386] = !f[406] && f[517] && f[212] && f[233]; // c3t943i94
	assign leaf[1387] = f[406] && !f[466] && !f[300] && !f[544]; // c3t943i94
	assign leaf[1388] = f[406] && !f[466] && !f[300] && f[544]; // c3t943i94
	assign leaf[1389] = f[406] && !f[466] && f[300] && !f[574]; // c3t943i94
	assign leaf[1390] = f[406] && !f[466] && f[300] && f[574]; // c3t943i94
	assign leaf[1391] = f[406] && f[466] && !f[347] && !f[291]; // c3t943i94
	assign leaf[1392] = f[406] && f[466] && !f[347] && f[291]; // c3t943i94
	assign leaf[1393] = f[406] && f[466] && f[347] && !f[318]; // c3t943i94
	assign leaf[1394] = f[406] && f[466] && f[347] && f[318]; // c3t943i94
	assign leaf[1395] = !f[401] && !f[347] && !f[321] && !f[570]; // c3t953i95
	assign leaf[1396] = !f[401] && !f[347] && !f[321] && f[570]; // c3t953i95
	assign leaf[1397] = !f[401] && !f[347] && f[321] && !f[127]; // c3t953i95
	assign leaf[1398] = !f[401] && !f[347] && f[321] && f[127]; // c3t953i95
	assign leaf[1399] = !f[401] && f[347] && !f[321] && !f[174]; // c3t953i95
	assign leaf[1400] = !f[401] && f[347] && !f[321] && f[174]; // c3t953i95
	assign leaf[1401] = !f[401] && f[347] && f[321] && !f[430]; // c3t953i95
	assign leaf[1402] = !f[401] && f[347] && f[321] && f[430]; // c3t953i95
	assign leaf[1403] = f[401] && !f[651] && !f[384] && !f[328]; // c3t953i95
	assign leaf[1404] = f[401] && !f[651] && !f[384] && f[328]; // c3t953i95
	assign leaf[1405] = f[401] && !f[651] && f[384] && !f[292]; // c3t953i95
	assign leaf[1406] = f[401] && !f[651] && f[384] && f[292]; // c3t953i95
	assign leaf[1407] = f[401] && f[651] && !f[565] && !f[568]; // c3t953i95
	assign leaf[1408] = f[401] && f[651] && !f[565] && f[568]; // c3t953i95
	assign leaf[1409] = f[401] && f[651] && f[565] && !f[455]; // c3t953i95
	assign leaf[1410] = f[401] && f[651] && f[565] && f[455]; // c3t953i95
	assign leaf[1411] = !f[427] && !f[241] && !f[719] && !f[518]; // c3t963i96
	assign leaf[1412] = !f[427] && !f[241] && !f[719] && f[518]; // c3t963i96
	assign leaf[1413] = !f[427] && !f[241] && f[719]; // c3t963i96
	assign leaf[1414] = !f[427] && f[241] && !f[303] && !f[184]; // c3t963i96
	assign leaf[1415] = !f[427] && f[241] && !f[303] && f[184]; // c3t963i96
	assign leaf[1416] = !f[427] && f[241] && f[303] && !f[235]; // c3t963i96
	assign leaf[1417] = !f[427] && f[241] && f[303] && f[235]; // c3t963i96
	assign leaf[1418] = f[427] && !f[437] && !f[236] && !f[327]; // c3t963i96
	assign leaf[1419] = f[427] && !f[437] && !f[236] && f[327]; // c3t963i96
	assign leaf[1420] = f[427] && !f[437] && f[236] && !f[215]; // c3t963i96
	assign leaf[1421] = f[427] && !f[437] && f[236] && f[215]; // c3t963i96
	assign leaf[1422] = f[427] && f[437] && !f[428]; // c3t963i96
	assign leaf[1423] = f[427] && f[437] && f[428] && !f[241]; // c3t963i96
	assign leaf[1424] = f[427] && f[437] && f[428] && f[241]; // c3t963i96
	assign leaf[1425] = !f[492] && !f[598] && !f[575] && !f[600]; // c3t973i97
	assign leaf[1426] = !f[492] && !f[598] && !f[575] && f[600]; // c3t973i97
	assign leaf[1427] = !f[492] && !f[598] && f[575] && !f[354]; // c3t973i97
	assign leaf[1428] = !f[492] && !f[598] && f[575] && f[354]; // c3t973i97
	assign leaf[1429] = !f[492] && f[598] && !f[629] && !f[495]; // c3t973i97
	assign leaf[1430] = !f[492] && f[598] && !f[629] && f[495]; // c3t973i97
	assign leaf[1431] = !f[492] && f[598] && f[629] && !f[573]; // c3t973i97
	assign leaf[1432] = !f[492] && f[598] && f[629] && f[573]; // c3t973i97
	assign leaf[1433] = f[492] && !f[468] && !f[493] && !f[293]; // c3t973i97
	assign leaf[1434] = f[492] && !f[468] && !f[493] && f[293]; // c3t973i97
	assign leaf[1435] = f[492] && !f[468] && f[493] && !f[346]; // c3t973i97
	assign leaf[1436] = f[492] && !f[468] && f[493] && f[346]; // c3t973i97
	assign leaf[1437] = f[492] && f[468] && !f[554] && !f[274]; // c3t973i97
	assign leaf[1438] = f[492] && f[468] && !f[554] && f[274]; // c3t973i97
	assign leaf[1439] = f[492] && f[468] && f[554] && !f[297]; // c3t973i97
	assign leaf[1440] = f[492] && f[468] && f[554] && f[297]; // c3t973i97
	assign leaf[1441] = !f[240] && !f[189] && !f[356] && !f[129]; // c3t983i98
	assign leaf[1442] = !f[240] && !f[189] && !f[356] && f[129]; // c3t983i98
	assign leaf[1443] = !f[240] && !f[189] && f[356] && !f[155]; // c3t983i98
	assign leaf[1444] = !f[240] && !f[189] && f[356] && f[155]; // c3t983i98
	assign leaf[1445] = !f[240] && f[189] && !f[245] && !f[237]; // c3t983i98
	assign leaf[1446] = !f[240] && f[189] && !f[245] && f[237]; // c3t983i98
	assign leaf[1447] = !f[240] && f[189] && f[245] && !f[627]; // c3t983i98
	assign leaf[1448] = !f[240] && f[189] && f[245] && f[627]; // c3t983i98
	assign leaf[1449] = f[240] && !f[128] && !f[319] && !f[209]; // c3t983i98
	assign leaf[1450] = f[240] && !f[128] && !f[319] && f[209]; // c3t983i98
	assign leaf[1451] = f[240] && !f[128] && f[319] && !f[316]; // c3t983i98
	assign leaf[1452] = f[240] && !f[128] && f[319] && f[316]; // c3t983i98
	assign leaf[1453] = f[240] && f[128] && !f[293] && !f[404]; // c3t983i98
	assign leaf[1454] = f[240] && f[128] && !f[293] && f[404]; // c3t983i98
	assign leaf[1455] = f[240] && f[128] && f[293] && !f[244]; // c3t983i98
	assign leaf[1456] = f[240] && f[128] && f[293] && f[244]; // c3t983i98
	assign leaf[1457] = !f[411] && !f[466] && !f[179] && !f[493]; // c3t993i99
	assign leaf[1458] = !f[411] && !f[466] && !f[179] && f[493]; // c3t993i99
	assign leaf[1459] = !f[411] && !f[466] && f[179] && !f[571]; // c3t993i99
	assign leaf[1460] = !f[411] && !f[466] && f[179] && f[571]; // c3t993i99
	assign leaf[1461] = !f[411] && f[466] && !f[382] && !f[548]; // c3t993i99
	assign leaf[1462] = !f[411] && f[466] && !f[382] && f[548]; // c3t993i99
	assign leaf[1463] = !f[411] && f[466] && f[382] && !f[356]; // c3t993i99
	assign leaf[1464] = !f[411] && f[466] && f[382] && f[356]; // c3t993i99
	assign leaf[1465] = f[411] && !f[179] && !f[235] && !f[130]; // c3t993i99
	assign leaf[1466] = f[411] && !f[179] && !f[235] && f[130]; // c3t993i99
	assign leaf[1467] = f[411] && !f[179] && f[235] && !f[464]; // c3t993i99
	assign leaf[1468] = f[411] && !f[179] && f[235] && f[464]; // c3t993i99
	assign leaf[1469] = f[411] && f[179] && !f[293] && !f[264]; // c3t993i99
	assign leaf[1470] = f[411] && f[179] && !f[293] && f[264]; // c3t993i99
	assign leaf[1471] = f[411] && f[179] && f[293] && !f[234]; // c3t993i99
	assign leaf[1472] = f[411] && f[179] && f[293] && f[234]; // c3t993i99
endmodule

module decision_tree_leaves_4(input logic [0:783] f, output logic [0:1315] leaf);
	assign leaf[0] = !f[211] && !f[428] && !f[402] && !f[398]; // c4t4i0
	assign leaf[1] = !f[211] && !f[428] && !f[402] && f[398]; // c4t4i0
	assign leaf[2] = !f[211] && !f[428] && f[402] && !f[155]; // c4t4i0
	assign leaf[3] = !f[211] && !f[428] && f[402] && f[155]; // c4t4i0
	assign leaf[4] = !f[211] && f[428] && !f[570] && !f[267]; // c4t4i0
	assign leaf[5] = !f[211] && f[428] && !f[570] && f[267]; // c4t4i0
	assign leaf[6] = !f[211] && f[428] && f[570] && !f[191]; // c4t4i0
	assign leaf[7] = !f[211] && f[428] && f[570] && f[191]; // c4t4i0
	assign leaf[8] = f[211] && !f[429] && !f[373] && !f[375]; // c4t4i0
	assign leaf[9] = f[211] && !f[429] && !f[373] && f[375]; // c4t4i0
	assign leaf[10] = f[211] && !f[429] && f[373] && !f[208]; // c4t4i0
	assign leaf[11] = f[211] && !f[429] && f[373] && f[208]; // c4t4i0
	assign leaf[12] = f[211] && f[429] && !f[210] && !f[600]; // c4t4i0
	assign leaf[13] = f[211] && f[429] && !f[210] && f[600]; // c4t4i0
	assign leaf[14] = f[211] && f[429] && f[210] && !f[213]; // c4t4i0
	assign leaf[15] = f[211] && f[429] && f[210] && f[213]; // c4t4i0
	assign leaf[16] = !f[400] && !f[402] && !f[398] && !f[375]; // c4t14i1
	assign leaf[17] = !f[400] && !f[402] && !f[398] && f[375]; // c4t14i1
	assign leaf[18] = !f[400] && !f[402] && f[398] && !f[458]; // c4t14i1
	assign leaf[19] = !f[400] && !f[402] && f[398] && f[458]; // c4t14i1
	assign leaf[20] = !f[400] && f[402] && !f[183] && !f[239]; // c4t14i1
	assign leaf[21] = !f[400] && f[402] && !f[183] && f[239]; // c4t14i1
	assign leaf[22] = !f[400] && f[402] && f[183] && !f[185]; // c4t14i1
	assign leaf[23] = !f[400] && f[402] && f[183] && f[185]; // c4t14i1
	assign leaf[24] = f[400] && !f[210] && !f[154] && !f[266]; // c4t14i1
	assign leaf[25] = f[400] && !f[210] && !f[154] && f[266]; // c4t14i1
	assign leaf[26] = f[400] && !f[210] && f[154] && !f[155]; // c4t14i1
	assign leaf[27] = f[400] && !f[210] && f[154] && f[155]; // c4t14i1
	assign leaf[28] = f[400] && f[210] && !f[463] && !f[628]; // c4t14i1
	assign leaf[29] = f[400] && f[210] && !f[463] && f[628]; // c4t14i1
	assign leaf[30] = f[400] && f[210] && f[463] && !f[212]; // c4t14i1
	assign leaf[31] = f[400] && f[210] && f[463] && f[212]; // c4t14i1
	assign leaf[32] = !f[183] && !f[267] && !f[437] && !f[464]; // c4t24i2
	assign leaf[33] = !f[183] && !f[267] && !f[437] && f[464]; // c4t24i2
	assign leaf[34] = !f[183] && !f[267] && f[437] && !f[126]; // c4t24i2
	assign leaf[35] = !f[183] && !f[267] && f[437] && f[126]; // c4t24i2
	assign leaf[36] = !f[183] && f[267] && !f[429] && !f[375]; // c4t24i2
	assign leaf[37] = !f[183] && f[267] && !f[429] && f[375]; // c4t24i2
	assign leaf[38] = !f[183] && f[267] && f[429] && !f[237]; // c4t24i2
	assign leaf[39] = !f[183] && f[267] && f[429] && f[237]; // c4t24i2
	assign leaf[40] = f[183] && !f[180] && !f[662] && !f[464]; // c4t24i2
	assign leaf[41] = f[183] && !f[180] && !f[662] && f[464]; // c4t24i2
	assign leaf[42] = f[183] && !f[180] && f[662] && !f[235]; // c4t24i2
	assign leaf[43] = f[183] && !f[180] && f[662] && f[235]; // c4t24i2
	assign leaf[44] = f[183] && f[180] && !f[182] && !f[153]; // c4t24i2
	assign leaf[45] = f[183] && f[180] && !f[182] && f[153]; // c4t24i2
	assign leaf[46] = f[183] && f[180] && f[182] && !f[184]; // c4t24i2
	assign leaf[47] = f[183] && f[180] && f[182] && f[184]; // c4t24i2
	assign leaf[48] = !f[401] && !f[399] && !f[374] && !f[397]; // c4t34i3
	assign leaf[49] = !f[401] && !f[399] && !f[374] && f[397]; // c4t34i3
	assign leaf[50] = !f[401] && !f[399] && f[374] && !f[184]; // c4t34i3
	assign leaf[51] = !f[401] && !f[399] && f[374] && f[184]; // c4t34i3
	assign leaf[52] = !f[401] && f[399] && !f[458] && !f[487]; // c4t34i3
	assign leaf[53] = !f[401] && f[399] && !f[458] && f[487]; // c4t34i3
	assign leaf[54] = !f[401] && f[399] && f[458] && !f[210]; // c4t34i3
	assign leaf[55] = !f[401] && f[399] && f[458] && f[210]; // c4t34i3
	assign leaf[56] = f[401] && !f[569] && !f[463] && !f[210]; // c4t34i3
	assign leaf[57] = f[401] && !f[569] && !f[463] && f[210]; // c4t34i3
	assign leaf[58] = f[401] && !f[569] && f[463] && !f[209]; // c4t34i3
	assign leaf[59] = f[401] && !f[569] && f[463] && f[209]; // c4t34i3
	assign leaf[60] = f[401] && f[569] && !f[488] && !f[136]; // c4t34i3
	assign leaf[61] = f[401] && f[569] && !f[488] && f[136]; // c4t34i3
	assign leaf[62] = f[401] && f[569] && f[488] && !f[574]; // c4t34i3
	assign leaf[63] = f[401] && f[569] && f[488] && f[574]; // c4t34i3
	assign leaf[64] = !f[597] && !f[210] && !f[543] && !f[266]; // c4t44i4
	assign leaf[65] = !f[597] && !f[210] && !f[543] && f[266]; // c4t44i4
	assign leaf[66] = !f[597] && !f[210] && f[543] && !f[189]; // c4t44i4
	assign leaf[67] = !f[597] && !f[210] && f[543] && f[189]; // c4t44i4
	assign leaf[68] = !f[597] && f[210] && !f[319] && !f[208]; // c4t44i4
	assign leaf[69] = !f[597] && f[210] && !f[319] && f[208]; // c4t44i4
	assign leaf[70] = !f[597] && f[210] && f[319] && !f[455]; // c4t44i4
	assign leaf[71] = !f[597] && f[210] && f[319] && f[455]; // c4t44i4
	assign leaf[72] = f[597] && !f[163] && !f[220] && !f[156]; // c4t44i4
	assign leaf[73] = f[597] && !f[163] && !f[220] && f[156]; // c4t44i4
	assign leaf[74] = f[597] && !f[163] && f[220] && !f[243]; // c4t44i4
	assign leaf[75] = f[597] && !f[163] && f[220] && f[243]; // c4t44i4
	assign leaf[76] = f[597] && f[163] && !f[187] && !f[567]; // c4t44i4
	assign leaf[77] = f[597] && f[163] && !f[187] && f[567]; // c4t44i4
	assign leaf[78] = f[597] && f[163] && f[187] && !f[213]; // c4t44i4
	assign leaf[79] = f[597] && f[163] && f[187] && f[213]; // c4t44i4
	assign leaf[80] = !f[464] && !f[183] && !f[436] && !f[295]; // c4t54i5
	assign leaf[81] = !f[464] && !f[183] && !f[436] && f[295]; // c4t54i5
	assign leaf[82] = !f[464] && !f[183] && f[436] && !f[575]; // c4t54i5
	assign leaf[83] = !f[464] && !f[183] && f[436] && f[575]; // c4t54i5
	assign leaf[84] = !f[464] && f[183] && !f[185] && !f[246]; // c4t54i5
	assign leaf[85] = !f[464] && f[183] && !f[185] && f[246]; // c4t54i5
	assign leaf[86] = !f[464] && f[183] && f[185] && !f[368]; // c4t54i5
	assign leaf[87] = !f[464] && f[183] && f[185] && f[368]; // c4t54i5
	assign leaf[88] = f[464] && !f[210] && !f[154] && !f[266]; // c4t54i5
	assign leaf[89] = f[464] && !f[210] && !f[154] && f[266]; // c4t54i5
	assign leaf[90] = f[464] && !f[210] && f[154] && !f[155]; // c4t54i5
	assign leaf[91] = f[464] && !f[210] && f[154] && f[155]; // c4t54i5
	assign leaf[92] = f[464] && f[210] && !f[213] && !f[292]; // c4t54i5
	assign leaf[93] = f[464] && f[210] && !f[213] && f[292]; // c4t54i5
	assign leaf[94] = f[464] && f[210] && f[213] && !f[442]; // c4t54i5
	assign leaf[95] = f[464] && f[210] && f[213] && f[442]; // c4t54i5
	assign leaf[96] = !f[569] && !f[427] && !f[374] && !f[373]; // c4t64i6
	assign leaf[97] = !f[569] && !f[427] && !f[374] && f[373]; // c4t64i6
	assign leaf[98] = !f[569] && !f[427] && f[374] && !f[551]; // c4t64i6
	assign leaf[99] = !f[569] && !f[427] && f[374] && f[551]; // c4t64i6
	assign leaf[100] = !f[569] && f[427] && !f[374] && !f[238]; // c4t64i6
	assign leaf[101] = !f[569] && f[427] && !f[374] && f[238]; // c4t64i6
	assign leaf[102] = !f[569] && f[427] && f[374] && !f[623]; // c4t64i6
	assign leaf[103] = !f[569] && f[427] && f[374] && f[623]; // c4t64i6
	assign leaf[104] = f[569] && !f[163] && !f[600] && !f[400]; // c4t64i6
	assign leaf[105] = f[569] && !f[163] && !f[600] && f[400]; // c4t64i6
	assign leaf[106] = f[569] && !f[163] && f[600] && !f[710]; // c4t64i6
	assign leaf[107] = f[569] && !f[163] && f[600] && f[710]; // c4t64i6
	assign leaf[108] = f[569] && f[163] && !f[595] && !f[213]; // c4t64i6
	assign leaf[109] = f[569] && f[163] && !f[595] && f[213]; // c4t64i6
	assign leaf[110] = f[569] && f[163] && f[595] && !f[567]; // c4t64i6
	assign leaf[111] = f[569] && f[163] && f[595] && f[567]; // c4t64i6
	assign leaf[112] = !f[401] && !f[598] && !f[238] && !f[182]; // c4t74i7
	assign leaf[113] = !f[401] && !f[598] && !f[238] && f[182]; // c4t74i7
	assign leaf[114] = !f[401] && !f[598] && f[238] && !f[430]; // c4t74i7
	assign leaf[115] = !f[401] && !f[598] && f[238] && f[430]; // c4t74i7
	assign leaf[116] = !f[401] && f[598] && !f[163] && !f[681]; // c4t74i7
	assign leaf[117] = !f[401] && f[598] && !f[163] && f[681]; // c4t74i7
	assign leaf[118] = !f[401] && f[598] && f[163] && !f[595]; // c4t74i7
	assign leaf[119] = !f[401] && f[598] && f[163] && f[595]; // c4t74i7
	assign leaf[120] = f[401] && !f[552] && !f[462] && !f[626]; // c4t74i7
	assign leaf[121] = f[401] && !f[552] && !f[462] && f[626]; // c4t74i7
	assign leaf[122] = f[401] && !f[552] && f[462] && !f[567]; // c4t74i7
	assign leaf[123] = f[401] && !f[552] && f[462] && f[567]; // c4t74i7
	assign leaf[124] = f[401] && f[552] && !f[664] && !f[454]; // c4t74i7
	assign leaf[125] = f[401] && f[552] && !f[664] && f[454]; // c4t74i7
	assign leaf[126] = f[401] && f[552] && f[664] && !f[209]; // c4t74i7
	assign leaf[127] = f[401] && f[552] && f[664] && f[209]; // c4t74i7
	assign leaf[128] = !f[568] && !f[455] && !f[238] && !f[182]; // c4t84i8
	assign leaf[129] = !f[568] && !f[455] && !f[238] && f[182]; // c4t84i8
	assign leaf[130] = !f[568] && !f[455] && f[238] && !f[240]; // c4t84i8
	assign leaf[131] = !f[568] && !f[455] && f[238] && f[240]; // c4t84i8
	assign leaf[132] = !f[568] && f[455] && !f[347] && !f[238]; // c4t84i8
	assign leaf[133] = !f[568] && f[455] && !f[347] && f[238]; // c4t84i8
	assign leaf[134] = !f[568] && f[455] && f[347] && !f[491]; // c4t84i8
	assign leaf[135] = !f[568] && f[455] && f[347] && f[491]; // c4t84i8
	assign leaf[136] = f[568] && !f[626] && !f[135] && !f[381]; // c4t84i8
	assign leaf[137] = f[568] && !f[626] && !f[135] && f[381]; // c4t84i8
	assign leaf[138] = f[568] && !f[626] && f[135] && !f[598]; // c4t84i8
	assign leaf[139] = f[568] && !f[626] && f[135] && f[598]; // c4t84i8
	assign leaf[140] = f[568] && f[626] && !f[426] && !f[136]; // c4t84i8
	assign leaf[141] = f[568] && f[626] && !f[426] && f[136]; // c4t84i8
	assign leaf[142] = f[568] && f[626] && f[426] && !f[462]; // c4t84i8
	assign leaf[143] = f[568] && f[626] && f[426] && f[462]; // c4t84i8
	assign leaf[144] = !f[464] && !f[603] && !f[295] && !f[659]; // c4t94i9
	assign leaf[145] = !f[464] && !f[603] && !f[295] && f[659]; // c4t94i9
	assign leaf[146] = !f[464] && !f[603] && f[295] && !f[346]; // c4t94i9
	assign leaf[147] = !f[464] && !f[603] && f[295] && f[346]; // c4t94i9
	assign leaf[148] = !f[464] && f[603] && !f[688] && !f[686]; // c4t94i9
	assign leaf[149] = !f[464] && f[603] && !f[688] && f[686]; // c4t94i9
	assign leaf[150] = !f[464] && f[603] && f[688] && !f[210]; // c4t94i9
	assign leaf[151] = !f[464] && f[603] && f[688] && f[210]; // c4t94i9
	assign leaf[152] = f[464] && !f[569] && !f[208] && !f[710]; // c4t94i9
	assign leaf[153] = f[464] && !f[569] && !f[208] && f[710]; // c4t94i9
	assign leaf[154] = f[464] && !f[569] && f[208] && !f[319]; // c4t94i9
	assign leaf[155] = f[464] && !f[569] && f[208] && f[319]; // c4t94i9
	assign leaf[156] = f[464] && f[569] && !f[163] && !f[399]; // c4t94i9
	assign leaf[157] = f[464] && f[569] && !f[163] && f[399]; // c4t94i9
	assign leaf[158] = f[464] && f[569] && f[163] && !f[213]; // c4t94i9
	assign leaf[159] = f[464] && f[569] && f[163] && f[213]; // c4t94i9
	assign leaf[160] = !f[463] && !f[628] && !f[322] && !f[238]; // c4t104i10
	assign leaf[161] = !f[463] && !f[628] && !f[322] && f[238]; // c4t104i10
	assign leaf[162] = !f[463] && !f[628] && f[322] && !f[375]; // c4t104i10
	assign leaf[163] = !f[463] && !f[628] && f[322] && f[375]; // c4t104i10
	assign leaf[164] = !f[463] && f[628] && !f[163] && !f[490]; // c4t104i10
	assign leaf[165] = !f[463] && f[628] && !f[163] && f[490]; // c4t104i10
	assign leaf[166] = !f[463] && f[628] && f[163] && !f[595]; // c4t104i10
	assign leaf[167] = !f[463] && f[628] && f[163] && f[595]; // c4t104i10
	assign leaf[168] = f[463] && !f[542] && !f[624] && !f[347]; // c4t104i10
	assign leaf[169] = f[463] && !f[542] && !f[624] && f[347]; // c4t104i10
	assign leaf[170] = f[463] && !f[542] && f[624] && !f[516]; // c4t104i10
	assign leaf[171] = f[463] && !f[542] && f[624] && f[516]; // c4t104i10
	assign leaf[172] = f[463] && f[542] && !f[163] && !f[220]; // c4t104i10
	assign leaf[173] = f[463] && f[542] && !f[163] && f[220]; // c4t104i10
	assign leaf[174] = f[463] && f[542] && f[163] && !f[213]; // c4t104i10
	assign leaf[175] = f[463] && f[542] && f[163] && f[213]; // c4t104i10
	assign leaf[176] = !f[437] && !f[577] && !f[322] && !f[239]; // c4t114i11
	assign leaf[177] = !f[437] && !f[577] && !f[322] && f[239]; // c4t114i11
	assign leaf[178] = !f[437] && !f[577] && f[322] && !f[408]; // c4t114i11
	assign leaf[179] = !f[437] && !f[577] && f[322] && f[408]; // c4t114i11
	assign leaf[180] = !f[437] && f[577] && !f[690] && !f[438]; // c4t114i11
	assign leaf[181] = !f[437] && f[577] && !f[690] && f[438]; // c4t114i11
	assign leaf[182] = !f[437] && f[577] && f[690] && !f[269]; // c4t114i11
	assign leaf[183] = !f[437] && f[577] && f[690] && f[269]; // c4t114i11
	assign leaf[184] = f[437] && !f[461] && !f[434] && !f[484]; // c4t114i11
	assign leaf[185] = f[437] && !f[461] && !f[434] && f[484]; // c4t114i11
	assign leaf[186] = f[437] && !f[461] && f[434] && !f[598]; // c4t114i11
	assign leaf[187] = f[437] && !f[461] && f[434] && f[598]; // c4t114i11
	assign leaf[188] = f[437] && f[461] && !f[542] && !f[234]; // c4t114i11
	assign leaf[189] = f[437] && f[461] && !f[542] && f[234]; // c4t114i11
	assign leaf[190] = f[437] && f[461] && f[542] && !f[183]; // c4t114i11
	assign leaf[191] = f[437] && f[461] && f[542] && f[183]; // c4t114i11
	assign leaf[192] = !f[346] && !f[208] && !f[465] && !f[637]; // c4t124i12
	assign leaf[193] = !f[346] && !f[208] && !f[465] && f[637]; // c4t124i12
	assign leaf[194] = !f[346] && !f[208] && f[465] && !f[291]; // c4t124i12
	assign leaf[195] = !f[346] && !f[208] && f[465] && f[291]; // c4t124i12
	assign leaf[196] = !f[346] && f[208] && !f[211] && !f[218]; // c4t124i12
	assign leaf[197] = !f[346] && f[208] && !f[211] && f[218]; // c4t124i12
	assign leaf[198] = !f[346] && f[208] && f[211] && !f[248]; // c4t124i12
	assign leaf[199] = !f[346] && f[208] && f[211] && f[248]; // c4t124i12
	assign leaf[200] = f[346] && !f[427] && !f[551] && !f[238]; // c4t124i12
	assign leaf[201] = f[346] && !f[427] && !f[551] && f[238]; // c4t124i12
	assign leaf[202] = f[346] && !f[427] && f[551] && !f[603]; // c4t124i12
	assign leaf[203] = f[346] && !f[427] && f[551] && f[603]; // c4t124i12
	assign leaf[204] = f[346] && f[427] && !f[568] && !f[710]; // c4t124i12
	assign leaf[205] = f[346] && f[427] && !f[568] && f[710]; // c4t124i12
	assign leaf[206] = f[346] && f[427] && f[568] && !f[157]; // c4t124i12
	assign leaf[207] = f[346] && f[427] && f[568] && f[157]; // c4t124i12
	assign leaf[208] = !f[595] && !f[374] && !f[426] && !f[373]; // c4t134i13
	assign leaf[209] = !f[595] && !f[374] && !f[426] && f[373]; // c4t134i13
	assign leaf[210] = !f[595] && !f[374] && f[426] && !f[294]; // c4t134i13
	assign leaf[211] = !f[595] && !f[374] && f[426] && f[294]; // c4t134i13
	assign leaf[212] = !f[595] && f[374] && !f[552] && !f[712]; // c4t134i13
	assign leaf[213] = !f[595] && f[374] && !f[552] && f[712]; // c4t134i13
	assign leaf[214] = !f[595] && f[374] && f[552] && !f[454]; // c4t134i13
	assign leaf[215] = !f[595] && f[374] && f[552] && f[454]; // c4t134i13
	assign leaf[216] = f[595] && !f[542] && !f[664]; // c4t134i13
	assign leaf[217] = f[595] && !f[542] && f[664]; // c4t134i13
	assign leaf[218] = f[595] && f[542] && !f[401] && !f[442]; // c4t134i13
	assign leaf[219] = f[595] && f[542] && !f[401] && f[442]; // c4t134i13
	assign leaf[220] = f[595] && f[542] && f[401] && !f[567]; // c4t134i13
	assign leaf[221] = f[595] && f[542] && f[401] && f[567]; // c4t134i13
	assign leaf[222] = !f[408] && !f[466] && !f[146] && !f[381]; // c4t144i14
	assign leaf[223] = !f[408] && !f[466] && !f[146] && f[381]; // c4t144i14
	assign leaf[224] = !f[408] && !f[466] && f[146]; // c4t144i14
	assign leaf[225] = !f[408] && f[466] && !f[488] && !f[295]; // c4t144i14
	assign leaf[226] = !f[408] && f[466] && !f[488] && f[295]; // c4t144i14
	assign leaf[227] = !f[408] && f[466] && f[488] && !f[572]; // c4t144i14
	assign leaf[228] = !f[408] && f[466] && f[488] && f[572]; // c4t144i14
	assign leaf[229] = f[408] && !f[209] && !f[544] && !f[627]; // c4t144i14
	assign leaf[230] = f[408] && !f[209] && !f[544] && f[627]; // c4t144i14
	assign leaf[231] = f[408] && !f[209] && f[544] && !f[551]; // c4t144i14
	assign leaf[232] = f[408] && !f[209] && f[544] && f[551]; // c4t144i14
	assign leaf[233] = f[408] && f[209] && !f[212] && !f[205]; // c4t144i14
	assign leaf[234] = f[408] && f[209] && !f[212] && f[205]; // c4t144i14
	assign leaf[235] = f[408] && f[209] && f[212] && !f[320]; // c4t144i14
	assign leaf[236] = f[408] && f[209] && f[212] && f[320]; // c4t144i14
	assign leaf[237] = !f[427] && !f[375] && !f[293] && !f[209]; // c4t154i15
	assign leaf[238] = !f[427] && !f[375] && !f[293] && f[209]; // c4t154i15
	assign leaf[239] = !f[427] && !f[375] && f[293] && !f[190]; // c4t154i15
	assign leaf[240] = !f[427] && !f[375] && f[293] && f[190]; // c4t154i15
	assign leaf[241] = !f[427] && f[375] && !f[408] && !f[409]; // c4t154i15
	assign leaf[242] = !f[427] && f[375] && !f[408] && f[409]; // c4t154i15
	assign leaf[243] = !f[427] && f[375] && f[408] && !f[601]; // c4t154i15
	assign leaf[244] = !f[427] && f[375] && f[408] && f[601]; // c4t154i15
	assign leaf[245] = f[427] && !f[346] && !f[237] && !f[181]; // c4t154i15
	assign leaf[246] = f[427] && !f[346] && !f[237] && f[181]; // c4t154i15
	assign leaf[247] = f[427] && !f[346] && f[237] && !f[191]; // c4t154i15
	assign leaf[248] = f[427] && !f[346] && f[237] && f[191]; // c4t154i15
	assign leaf[249] = f[427] && f[346] && !f[328] && !f[325]; // c4t154i15
	assign leaf[250] = f[427] && f[346] && !f[328] && f[325]; // c4t154i15
	assign leaf[251] = f[427] && f[346] && f[328] && !f[241]; // c4t154i15
	assign leaf[252] = f[427] && f[346] && f[328] && f[241]; // c4t154i15
	assign leaf[253] = !f[568] && !f[454] && !f[375] && !f[401]; // c4t164i16
	assign leaf[254] = !f[568] && !f[454] && !f[375] && f[401]; // c4t164i16
	assign leaf[255] = !f[568] && !f[454] && f[375] && !f[551]; // c4t164i16
	assign leaf[256] = !f[568] && !f[454] && f[375] && f[551]; // c4t164i16
	assign leaf[257] = !f[568] && f[454] && !f[331] && !f[345]; // c4t164i16
	assign leaf[258] = !f[568] && f[454] && !f[331] && f[345]; // c4t164i16
	assign leaf[259] = !f[568] && f[454] && f[331] && !f[209]; // c4t164i16
	assign leaf[260] = !f[568] && f[454] && f[331] && f[209]; // c4t164i16
	assign leaf[261] = f[568] && !f[626] && !f[636] && !f[298]; // c4t164i16
	assign leaf[262] = f[568] && !f[626] && !f[636] && f[298]; // c4t164i16
	assign leaf[263] = f[568] && !f[626] && f[636] && !f[182]; // c4t164i16
	assign leaf[264] = f[568] && !f[626] && f[636] && f[182]; // c4t164i16
	assign leaf[265] = f[568] && f[626] && !f[399]; // c4t164i16
	assign leaf[266] = f[568] && f[626] && f[399] && !f[628]; // c4t164i16
	assign leaf[267] = f[568] && f[626] && f[399] && f[628]; // c4t164i16
	assign leaf[268] = !f[463] && !f[628] && !f[323] && !f[574]; // c4t174i17
	assign leaf[269] = !f[463] && !f[628] && !f[323] && f[574]; // c4t174i17
	assign leaf[270] = !f[463] && !f[628] && f[323] && !f[380]; // c4t174i17
	assign leaf[271] = !f[463] && !f[628] && f[323] && f[380]; // c4t174i17
	assign leaf[272] = !f[463] && f[628] && !f[462] && !f[219]; // c4t174i17
	assign leaf[273] = !f[463] && f[628] && !f[462] && f[219]; // c4t174i17
	assign leaf[274] = !f[463] && f[628] && f[462] && !f[347]; // c4t174i17
	assign leaf[275] = !f[463] && f[628] && f[462] && f[347]; // c4t174i17
	assign leaf[276] = f[463] && !f[740] && !f[542] && !f[208]; // c4t174i17
	assign leaf[277] = f[463] && !f[740] && !f[542] && f[208]; // c4t174i17
	assign leaf[278] = f[463] && !f[740] && f[542] && !f[163]; // c4t174i17
	assign leaf[279] = f[463] && !f[740] && f[542] && f[163]; // c4t174i17
	assign leaf[280] = f[463] && f[740] && !f[426]; // c4t174i17
	assign leaf[281] = f[463] && f[740] && f[426]; // c4t174i17
	assign leaf[282] = !f[594] && !f[208] && !f[601] && !f[657]; // c4t184i18
	assign leaf[283] = !f[594] && !f[208] && !f[601] && f[657]; // c4t184i18
	assign leaf[284] = !f[594] && !f[208] && f[601] && !f[490]; // c4t184i18
	assign leaf[285] = !f[594] && !f[208] && f[601] && f[490]; // c4t184i18
	assign leaf[286] = !f[594] && f[208] && !f[184] && !f[239]; // c4t184i18
	assign leaf[287] = !f[594] && f[208] && !f[184] && f[239]; // c4t184i18
	assign leaf[288] = !f[594] && f[208] && f[184] && !f[183]; // c4t184i18
	assign leaf[289] = !f[594] && f[208] && f[184] && f[183]; // c4t184i18
	assign leaf[290] = f[594] && !f[527] && !f[372]; // c4t184i18
	assign leaf[291] = f[594] && !f[527] && f[372] && !f[625]; // c4t184i18
	assign leaf[292] = f[594] && !f[527] && f[372] && f[625]; // c4t184i18
	assign leaf[293] = f[594] && f[527]; // c4t184i18
	assign leaf[294] = !f[491] && !f[629] && !f[236] && !f[180]; // c4t194i19
	assign leaf[295] = !f[491] && !f[629] && !f[236] && f[180]; // c4t194i19
	assign leaf[296] = !f[491] && !f[629] && f[236] && !f[291]; // c4t194i19
	assign leaf[297] = !f[491] && !f[629] && f[236] && f[291]; // c4t194i19
	assign leaf[298] = !f[491] && f[629] && !f[630] && !f[490]; // c4t194i19
	assign leaf[299] = !f[491] && f[629] && !f[630] && f[490]; // c4t194i19
	assign leaf[300] = !f[491] && f[629] && f[630] && !f[302]; // c4t194i19
	assign leaf[301] = !f[491] && f[629] && f[630] && f[302]; // c4t194i19
	assign leaf[302] = f[491] && !f[466] && !f[212] && !f[295]; // c4t194i19
	assign leaf[303] = f[491] && !f[466] && !f[212] && f[295]; // c4t194i19
	assign leaf[304] = f[491] && !f[466] && f[212] && !f[296]; // c4t194i19
	assign leaf[305] = f[491] && !f[466] && f[212] && f[296]; // c4t194i19
	assign leaf[306] = f[491] && f[466] && !f[260] && !f[383]; // c4t194i19
	assign leaf[307] = f[491] && f[466] && !f[260] && f[383]; // c4t194i19
	assign leaf[308] = f[491] && f[466] && f[260] && !f[293]; // c4t194i19
	assign leaf[309] = f[491] && f[466] && f[260] && f[293]; // c4t194i19
	assign leaf[310] = !f[409] && !f[405] && !f[488] && !f[460]; // c4t204i20
	assign leaf[311] = !f[409] && !f[405] && !f[488] && f[460]; // c4t204i20
	assign leaf[312] = !f[409] && !f[405] && f[488] && !f[490]; // c4t204i20
	assign leaf[313] = !f[409] && !f[405] && f[488] && f[490]; // c4t204i20
	assign leaf[314] = !f[409] && f[405] && !f[521] && !f[346]; // c4t204i20
	assign leaf[315] = !f[409] && f[405] && !f[521] && f[346]; // c4t204i20
	assign leaf[316] = !f[409] && f[405] && f[521] && !f[410]; // c4t204i20
	assign leaf[317] = !f[409] && f[405] && f[521] && f[410]; // c4t204i20
	assign leaf[318] = f[409] && !f[375] && !f[265] && !f[182]; // c4t204i20
	assign leaf[319] = f[409] && !f[375] && !f[265] && f[182]; // c4t204i20
	assign leaf[320] = f[409] && !f[375] && f[265] && !f[426]; // c4t204i20
	assign leaf[321] = f[409] && !f[375] && f[265] && f[426]; // c4t204i20
	assign leaf[322] = f[409] && f[375] && !f[213] && !f[296]; // c4t204i20
	assign leaf[323] = f[409] && f[375] && !f[213] && f[296]; // c4t204i20
	assign leaf[324] = f[409] && f[375] && f[213] && !f[296]; // c4t204i20
	assign leaf[325] = f[409] && f[375] && f[213] && f[296]; // c4t204i20
	assign leaf[326] = !f[491] && !f[629] && !f[322] && !f[657]; // c4t214i21
	assign leaf[327] = !f[491] && !f[629] && !f[322] && f[657]; // c4t214i21
	assign leaf[328] = !f[491] && !f[629] && f[322] && !f[289]; // c4t214i21
	assign leaf[329] = !f[491] && !f[629] && f[322] && f[289]; // c4t214i21
	assign leaf[330] = !f[491] && f[629] && !f[184] && !f[685]; // c4t214i21
	assign leaf[331] = !f[491] && f[629] && !f[184] && f[685]; // c4t214i21
	assign leaf[332] = !f[491] && f[629] && f[184]; // c4t214i21
	assign leaf[333] = f[491] && !f[214] && !f[269] && !f[551]; // c4t214i21
	assign leaf[334] = f[491] && !f[214] && !f[269] && f[551]; // c4t214i21
	assign leaf[335] = f[491] && !f[214] && f[269] && !f[270]; // c4t214i21
	assign leaf[336] = f[491] && !f[214] && f[269] && f[270]; // c4t214i21
	assign leaf[337] = f[491] && f[214] && !f[297] && !f[468]; // c4t214i21
	assign leaf[338] = f[491] && f[214] && !f[297] && f[468]; // c4t214i21
	assign leaf[339] = f[491] && f[214] && f[297] && !f[183]; // c4t214i21
	assign leaf[340] = f[491] && f[214] && f[297] && f[183]; // c4t214i21
	assign leaf[341] = !f[430] && !f[625] && !f[482] && !f[347]; // c4t224i22
	assign leaf[342] = !f[430] && !f[625] && !f[482] && f[347]; // c4t224i22
	assign leaf[343] = !f[430] && !f[625] && f[482] && !f[406]; // c4t224i22
	assign leaf[344] = !f[430] && !f[625] && f[482] && f[406]; // c4t224i22
	assign leaf[345] = !f[430] && f[625] && !f[406] && !f[458]; // c4t224i22
	assign leaf[346] = !f[430] && f[625] && !f[406] && f[458]; // c4t224i22
	assign leaf[347] = !f[430] && f[625] && f[406] && !f[186]; // c4t224i22
	assign leaf[348] = !f[430] && f[625] && f[406] && f[186]; // c4t224i22
	assign leaf[349] = f[430] && !f[552] && !f[462] && !f[629]; // c4t224i22
	assign leaf[350] = f[430] && !f[552] && !f[462] && f[629]; // c4t224i22
	assign leaf[351] = f[430] && !f[552] && f[462] && !f[214]; // c4t224i22
	assign leaf[352] = f[430] && !f[552] && f[462] && f[214]; // c4t224i22
	assign leaf[353] = f[430] && f[552] && !f[270] && !f[273]; // c4t224i22
	assign leaf[354] = f[430] && f[552] && !f[270] && f[273]; // c4t224i22
	assign leaf[355] = f[430] && f[552] && f[270] && !f[209]; // c4t224i22
	assign leaf[356] = f[430] && f[552] && f[270] && f[209]; // c4t224i22
	assign leaf[357] = !f[465] && !f[577] && !f[212] && !f[295]; // c4t234i23
	assign leaf[358] = !f[465] && !f[577] && !f[212] && f[295]; // c4t234i23
	assign leaf[359] = !f[465] && !f[577] && f[212] && !f[237]; // c4t234i23
	assign leaf[360] = !f[465] && !f[577] && f[212] && f[237]; // c4t234i23
	assign leaf[361] = !f[465] && f[577] && !f[662] && !f[688]; // c4t234i23
	assign leaf[362] = !f[465] && f[577] && !f[662] && f[688]; // c4t234i23
	assign leaf[363] = !f[465] && f[577] && f[662] && !f[179]; // c4t234i23
	assign leaf[364] = !f[465] && f[577] && f[662] && f[179]; // c4t234i23
	assign leaf[365] = f[465] && !f[235] && !f[179] && !f[571]; // c4t234i23
	assign leaf[366] = f[465] && !f[235] && !f[179] && f[571]; // c4t234i23
	assign leaf[367] = f[465] && !f[235] && f[179] && !f[262]; // c4t234i23
	assign leaf[368] = f[465] && !f[235] && f[179] && f[262]; // c4t234i23
	assign leaf[369] = f[465] && f[235] && !f[232] && !f[184]; // c4t234i23
	assign leaf[370] = f[465] && f[235] && !f[232] && f[184]; // c4t234i23
	assign leaf[371] = f[465] && f[235] && f[232] && !f[219]; // c4t234i23
	assign leaf[372] = f[465] && f[235] && f[232] && f[219]; // c4t234i23
	assign leaf[373] = !f[347] && !f[345] && !f[343] && !f[348]; // c4t244i24
	assign leaf[374] = !f[347] && !f[345] && !f[343] && f[348]; // c4t244i24
	assign leaf[375] = !f[347] && !f[345] && f[343] && !f[180]; // c4t244i24
	assign leaf[376] = !f[347] && !f[345] && f[343] && f[180]; // c4t244i24
	assign leaf[377] = !f[347] && f[345] && !f[454] && !f[236]; // c4t244i24
	assign leaf[378] = !f[347] && f[345] && !f[454] && f[236]; // c4t244i24
	assign leaf[379] = !f[347] && f[345] && f[454] && !f[320]; // c4t244i24
	assign leaf[380] = !f[347] && f[345] && f[454] && f[320]; // c4t244i24
	assign leaf[381] = f[347] && !f[408] && !f[324] && !f[382]; // c4t244i24
	assign leaf[382] = f[347] && !f[408] && !f[324] && f[382]; // c4t244i24
	assign leaf[383] = f[347] && !f[408] && f[324] && !f[407]; // c4t244i24
	assign leaf[384] = f[347] && !f[408] && f[324] && f[407]; // c4t244i24
	assign leaf[385] = f[347] && f[408] && !f[241] && !f[186]; // c4t244i24
	assign leaf[386] = f[347] && f[408] && !f[241] && f[186]; // c4t244i24
	assign leaf[387] = f[347] && f[408] && f[241] && !f[244]; // c4t244i24
	assign leaf[388] = f[347] && f[408] && f[241] && f[244]; // c4t244i24
	assign leaf[389] = !f[346] && !f[207] && !f[263] && !f[571]; // c4t254i25
	assign leaf[390] = !f[346] && !f[207] && !f[263] && f[571]; // c4t254i25
	assign leaf[391] = !f[346] && !f[207] && f[263] && !f[260]; // c4t254i25
	assign leaf[392] = !f[346] && !f[207] && f[263] && f[260]; // c4t254i25
	assign leaf[393] = !f[346] && f[207] && !f[290] && !f[319]; // c4t254i25
	assign leaf[394] = !f[346] && f[207] && !f[290] && f[319]; // c4t254i25
	assign leaf[395] = !f[346] && f[207] && f[290] && !f[183]; // c4t254i25
	assign leaf[396] = !f[346] && f[207] && f[290] && f[183]; // c4t254i25
	assign leaf[397] = f[346] && !f[428] && !f[572] && !f[627]; // c4t254i25
	assign leaf[398] = f[346] && !f[428] && !f[572] && f[627]; // c4t254i25
	assign leaf[399] = f[346] && !f[428] && f[572] && !f[575]; // c4t254i25
	assign leaf[400] = f[346] && !f[428] && f[572] && f[575]; // c4t254i25
	assign leaf[401] = f[346] && f[428] && !f[214] && !f[211]; // c4t254i25
	assign leaf[402] = f[346] && f[428] && !f[214] && f[211]; // c4t254i25
	assign leaf[403] = f[346] && f[428] && f[214] && !f[273]; // c4t254i25
	assign leaf[404] = f[346] && f[428] && f[214] && f[273]; // c4t254i25
	assign leaf[405] = !f[740] && !f[409] && !f[438] && !f[577]; // c4t264i26
	assign leaf[406] = !f[740] && !f[409] && !f[438] && f[577]; // c4t264i26
	assign leaf[407] = !f[740] && !f[409] && f[438] && !f[248]; // c4t264i26
	assign leaf[408] = !f[740] && !f[409] && f[438] && f[248]; // c4t264i26
	assign leaf[409] = !f[740] && f[409] && !f[403] && !f[454]; // c4t264i26
	assign leaf[410] = !f[740] && f[409] && !f[403] && f[454]; // c4t264i26
	assign leaf[411] = !f[740] && f[409] && f[403] && !f[434]; // c4t264i26
	assign leaf[412] = !f[740] && f[409] && f[403] && f[434]; // c4t264i26
	assign leaf[413] = f[740] && !f[412]; // c4t264i26
	assign leaf[414] = f[740] && f[412]; // c4t264i26
	assign leaf[415] = !f[743] && !f[96] && !f[628] && !f[684]; // c4t274i27
	assign leaf[416] = !f[743] && !f[96] && !f[628] && f[684]; // c4t274i27
	assign leaf[417] = !f[743] && !f[96] && f[628] && !f[604]; // c4t274i27
	assign leaf[418] = !f[743] && !f[96] && f[628] && f[604]; // c4t274i27
	assign leaf[419] = !f[743] && f[96] && !f[574]; // c4t274i27
	assign leaf[420] = !f[743] && f[96] && f[574]; // c4t274i27
	assign leaf[421] = f[743] && !f[459] && !f[295]; // c4t274i27
	assign leaf[422] = f[743] && !f[459] && f[295]; // c4t274i27
	assign leaf[423] = f[743] && f[459]; // c4t274i27
	assign leaf[424] = !f[491] && !f[630] && !f[744] && !f[526]; // c4t284i28
	assign leaf[425] = !f[491] && !f[630] && !f[744] && f[526]; // c4t284i28
	assign leaf[426] = !f[491] && !f[630] && f[744]; // c4t284i28
	assign leaf[427] = !f[491] && f[630] && !f[328] && !f[455]; // c4t284i28
	assign leaf[428] = !f[491] && f[630] && !f[328] && f[455]; // c4t284i28
	assign leaf[429] = !f[491] && f[630] && f[328] && !f[213]; // c4t284i28
	assign leaf[430] = !f[491] && f[630] && f[328] && f[213]; // c4t284i28
	assign leaf[431] = f[491] && !f[571] && !f[626] && !f[739]; // c4t284i28
	assign leaf[432] = f[491] && !f[571] && !f[626] && f[739]; // c4t284i28
	assign leaf[433] = f[491] && !f[571] && f[626] && !f[544]; // c4t284i28
	assign leaf[434] = f[491] && !f[571] && f[626] && f[544]; // c4t284i28
	assign leaf[435] = f[491] && f[571] && !f[186] && !f[654]; // c4t284i28
	assign leaf[436] = f[491] && f[571] && !f[186] && f[654]; // c4t284i28
	assign leaf[437] = f[491] && f[571] && f[186] && !f[497]; // c4t284i28
	assign leaf[438] = f[491] && f[571] && f[186] && f[497]; // c4t284i28
	assign leaf[439] = !f[286] && !f[594] && !f[348] && !f[345]; // c4t294i29
	assign leaf[440] = !f[286] && !f[594] && !f[348] && f[345]; // c4t294i29
	assign leaf[441] = !f[286] && !f[594] && f[348] && !f[381]; // c4t294i29
	assign leaf[442] = !f[286] && !f[594] && f[348] && f[381]; // c4t294i29
	assign leaf[443] = !f[286] && f[594] && !f[553] && !f[206]; // c4t294i29
	assign leaf[444] = !f[286] && f[594] && !f[553] && f[206]; // c4t294i29
	assign leaf[445] = !f[286] && f[594] && f[553]; // c4t294i29
	assign leaf[446] = f[286] && !f[262] && !f[207] && !f[471]; // c4t294i29
	assign leaf[447] = f[286] && !f[262] && !f[207] && f[471]; // c4t294i29
	assign leaf[448] = f[286] && !f[262] && f[207] && !f[381]; // c4t294i29
	assign leaf[449] = f[286] && !f[262] && f[207] && f[381]; // c4t294i29
	assign leaf[450] = f[286] && f[262] && !f[218] && !f[396]; // c4t294i29
	assign leaf[451] = f[286] && f[262] && !f[218] && f[396]; // c4t294i29
	assign leaf[452] = f[286] && f[262] && f[218] && !f[412]; // c4t294i29
	assign leaf[453] = f[286] && f[262] && f[218] && f[412]; // c4t294i29
	assign leaf[454] = !f[745] && !f[399] && !f[375] && !f[373]; // c4t304i30
	assign leaf[455] = !f[745] && !f[399] && !f[375] && f[373]; // c4t304i30
	assign leaf[456] = !f[745] && !f[399] && f[375] && !f[601]; // c4t304i30
	assign leaf[457] = !f[745] && !f[399] && f[375] && f[601]; // c4t304i30
	assign leaf[458] = !f[745] && f[399] && !f[514] && !f[322]; // c4t304i30
	assign leaf[459] = !f[745] && f[399] && !f[514] && f[322]; // c4t304i30
	assign leaf[460] = !f[745] && f[399] && f[514] && !f[434]; // c4t304i30
	assign leaf[461] = !f[745] && f[399] && f[514] && f[434]; // c4t304i30
	assign leaf[462] = f[745] && !f[483]; // c4t304i30
	assign leaf[463] = f[745] && f[483]; // c4t304i30
	assign leaf[464] = !f[208] && !f[327] && !f[352] && !f[272]; // c4t314i31
	assign leaf[465] = !f[208] && !f[327] && !f[352] && f[272]; // c4t314i31
	assign leaf[466] = !f[208] && !f[327] && f[352] && !f[436]; // c4t314i31
	assign leaf[467] = !f[208] && !f[327] && f[352] && f[436]; // c4t314i31
	assign leaf[468] = !f[208] && f[327] && !f[241] && !f[296]; // c4t314i31
	assign leaf[469] = !f[208] && f[327] && !f[241] && f[296]; // c4t314i31
	assign leaf[470] = !f[208] && f[327] && f[241] && !f[467]; // c4t314i31
	assign leaf[471] = !f[208] && f[327] && f[241] && f[467]; // c4t314i31
	assign leaf[472] = f[208] && !f[184] && !f[239] && !f[243]; // c4t314i31
	assign leaf[473] = f[208] && !f[184] && !f[239] && f[243]; // c4t314i31
	assign leaf[474] = f[208] && !f[184] && f[239] && !f[234]; // c4t314i31
	assign leaf[475] = f[208] && !f[184] && f[239] && f[234]; // c4t314i31
	assign leaf[476] = f[208] && f[184] && !f[182] && !f[296]; // c4t314i31
	assign leaf[477] = f[208] && f[184] && !f[182] && f[296]; // c4t314i31
	assign leaf[478] = f[208] && f[184] && f[182] && !f[248]; // c4t314i31
	assign leaf[479] = f[208] && f[184] && f[182] && f[248]; // c4t314i31
	assign leaf[480] = !f[219] && !f[286] && !f[600] && !f[655]; // c4t324i32
	assign leaf[481] = !f[219] && !f[286] && !f[600] && f[655]; // c4t324i32
	assign leaf[482] = !f[219] && !f[286] && f[600] && !f[576]; // c4t324i32
	assign leaf[483] = !f[219] && !f[286] && f[600] && f[576]; // c4t324i32
	assign leaf[484] = !f[219] && f[286] && !f[234] && !f[290]; // c4t324i32
	assign leaf[485] = !f[219] && f[286] && !f[234] && f[290]; // c4t324i32
	assign leaf[486] = !f[219] && f[286] && f[234] && !f[329]; // c4t324i32
	assign leaf[487] = !f[219] && f[286] && f[234] && f[329]; // c4t324i32
	assign leaf[488] = f[219] && !f[242] && !f[323] && !f[187]; // c4t324i32
	assign leaf[489] = f[219] && !f[242] && !f[323] && f[187]; // c4t324i32
	assign leaf[490] = f[219] && !f[242] && f[323] && !f[487]; // c4t324i32
	assign leaf[491] = f[219] && !f[242] && f[323] && f[487]; // c4t324i32
	assign leaf[492] = f[219] && f[242] && !f[240] && !f[655]; // c4t324i32
	assign leaf[493] = f[219] && f[242] && !f[240] && f[655]; // c4t324i32
	assign leaf[494] = f[219] && f[242] && f[240]; // c4t324i32
	assign leaf[495] = !f[490] && !f[411] && !f[236] && !f[268]; // c4t334i33
	assign leaf[496] = !f[490] && !f[411] && !f[236] && f[268]; // c4t334i33
	assign leaf[497] = !f[490] && !f[411] && f[236] && !f[262]; // c4t334i33
	assign leaf[498] = !f[490] && !f[411] && f[236] && f[262]; // c4t334i33
	assign leaf[499] = !f[490] && f[411] && !f[323] && !f[397]; // c4t334i33
	assign leaf[500] = !f[490] && f[411] && !f[323] && f[397]; // c4t334i33
	assign leaf[501] = !f[490] && f[411] && f[323] && !f[435]; // c4t334i33
	assign leaf[502] = !f[490] && f[411] && f[323] && f[435]; // c4t334i33
	assign leaf[503] = f[490] && !f[348] && !f[346] && !f[344]; // c4t334i33
	assign leaf[504] = f[490] && !f[348] && !f[346] && f[344]; // c4t334i33
	assign leaf[505] = f[490] && !f[348] && f[346] && !f[243]; // c4t334i33
	assign leaf[506] = f[490] && !f[348] && f[346] && f[243]; // c4t334i33
	assign leaf[507] = f[490] && f[348] && !f[322] && !f[186]; // c4t334i33
	assign leaf[508] = f[490] && f[348] && !f[322] && f[186]; // c4t334i33
	assign leaf[509] = f[490] && f[348] && f[322] && !f[211]; // c4t334i33
	assign leaf[510] = f[490] && f[348] && f[322] && f[211]; // c4t334i33
	assign leaf[511] = !f[746] && !f[456] && !f[408] && !f[322]; // c4t344i34
	assign leaf[512] = !f[746] && !f[456] && !f[408] && f[322]; // c4t344i34
	assign leaf[513] = !f[746] && !f[456] && f[408] && !f[524]; // c4t344i34
	assign leaf[514] = !f[746] && !f[456] && f[408] && f[524]; // c4t344i34
	assign leaf[515] = !f[746] && f[456] && !f[439] && !f[494]; // c4t344i34
	assign leaf[516] = !f[746] && f[456] && !f[439] && f[494]; // c4t344i34
	assign leaf[517] = !f[746] && f[456] && f[439] && !f[513]; // c4t344i34
	assign leaf[518] = !f[746] && f[456] && f[439] && f[513]; // c4t344i34
	assign leaf[519] = f[746]; // c4t344i34
	assign leaf[520] = !f[740] && !f[185] && !f[183] && !f[294]; // c4t354i35
	assign leaf[521] = !f[740] && !f[185] && !f[183] && f[294]; // c4t354i35
	assign leaf[522] = !f[740] && !f[185] && f[183] && !f[180]; // c4t354i35
	assign leaf[523] = !f[740] && !f[185] && f[183] && f[180]; // c4t354i35
	assign leaf[524] = !f[740] && f[185] && !f[296] && !f[294]; // c4t354i35
	assign leaf[525] = !f[740] && f[185] && !f[296] && f[294]; // c4t354i35
	assign leaf[526] = !f[740] && f[185] && f[296] && !f[182]; // c4t354i35
	assign leaf[527] = !f[740] && f[185] && f[296] && f[182]; // c4t354i35
	assign leaf[528] = f[740] && !f[240]; // c4t354i35
	assign leaf[529] = f[740] && f[240]; // c4t354i35
	assign leaf[530] = !f[744] && !f[128] && !f[739] && !f[747]; // c4t364i36
	assign leaf[531] = !f[744] && !f[128] && !f[739] && f[747]; // c4t364i36
	assign leaf[532] = !f[744] && !f[128] && f[739] && !f[412]; // c4t364i36
	assign leaf[533] = !f[744] && !f[128] && f[739] && f[412]; // c4t364i36
	assign leaf[534] = !f[744] && f[128] && !f[239] && !f[433]; // c4t364i36
	assign leaf[535] = !f[744] && f[128] && !f[239] && f[433]; // c4t364i36
	assign leaf[536] = !f[744] && f[128] && f[239] && !f[628]; // c4t364i36
	assign leaf[537] = !f[744] && f[128] && f[239] && f[628]; // c4t364i36
	assign leaf[538] = f[744] && !f[455] && !f[411]; // c4t364i36
	assign leaf[539] = f[744] && !f[455] && f[411]; // c4t364i36
	assign leaf[540] = f[744] && f[455]; // c4t364i36
	assign leaf[541] = !f[737] && !f[743] && !f[180] && !f[236]; // c4t374i37
	assign leaf[542] = !f[737] && !f[743] && !f[180] && f[236]; // c4t374i37
	assign leaf[543] = !f[737] && !f[743] && f[180] && !f[183]; // c4t374i37
	assign leaf[544] = !f[737] && !f[743] && f[180] && f[183]; // c4t374i37
	assign leaf[545] = !f[737] && f[743] && !f[298] && !f[353]; // c4t374i37
	assign leaf[546] = !f[737] && f[743] && !f[298] && f[353]; // c4t374i37
	assign leaf[547] = !f[737] && f[743] && f[298] && !f[490]; // c4t374i37
	assign leaf[548] = !f[737] && f[743] && f[298] && f[490]; // c4t374i37
	assign leaf[549] = f[737] && !f[385]; // c4t374i37
	assign leaf[550] = f[737] && f[385]; // c4t374i37
	assign leaf[551] = !f[332] && !f[737] && !f[185] && !f[187]; // c4t384i38
	assign leaf[552] = !f[332] && !f[737] && !f[185] && f[187]; // c4t384i38
	assign leaf[553] = !f[332] && !f[737] && f[185] && !f[182]; // c4t384i38
	assign leaf[554] = !f[332] && !f[737] && f[185] && f[182]; // c4t384i38
	assign leaf[555] = !f[332] && f[737] && !f[267]; // c4t384i38
	assign leaf[556] = !f[332] && f[737] && f[267]; // c4t384i38
	assign leaf[557] = f[332] && !f[371]; // c4t384i38
	assign leaf[558] = f[332] && f[371]; // c4t384i38
	assign leaf[559] = !f[96] && !f[409] && !f[405] && !f[516]; // c4t394i39
	assign leaf[560] = !f[96] && !f[409] && !f[405] && f[516]; // c4t394i39
	assign leaf[561] = !f[96] && !f[409] && f[405] && !f[326]; // c4t394i39
	assign leaf[562] = !f[96] && !f[409] && f[405] && f[326]; // c4t394i39
	assign leaf[563] = !f[96] && f[409] && !f[375] && !f[293]; // c4t394i39
	assign leaf[564] = !f[96] && f[409] && !f[375] && f[293]; // c4t394i39
	assign leaf[565] = !f[96] && f[409] && f[375] && !f[241]; // c4t394i39
	assign leaf[566] = !f[96] && f[409] && f[375] && f[241]; // c4t394i39
	assign leaf[567] = f[96] && !f[574]; // c4t394i39
	assign leaf[568] = f[96] && f[574]; // c4t394i39
	assign leaf[569] = !f[465] && !f[605] && !f[238] && !f[294]; // c4t404i40
	assign leaf[570] = !f[465] && !f[605] && !f[238] && f[294]; // c4t404i40
	assign leaf[571] = !f[465] && !f[605] && f[238] && !f[240]; // c4t404i40
	assign leaf[572] = !f[465] && !f[605] && f[238] && f[240]; // c4t404i40
	assign leaf[573] = !f[465] && f[605] && !f[218] && !f[662]; // c4t404i40
	assign leaf[574] = !f[465] && f[605] && !f[218] && f[662]; // c4t404i40
	assign leaf[575] = !f[465] && f[605] && f[218] && !f[291]; // c4t404i40
	assign leaf[576] = !f[465] && f[605] && f[218] && f[291]; // c4t404i40
	assign leaf[577] = f[465] && !f[381] && !f[297] && !f[214]; // c4t404i40
	assign leaf[578] = f[465] && !f[381] && !f[297] && f[214]; // c4t404i40
	assign leaf[579] = f[465] && !f[381] && f[297] && !f[549]; // c4t404i40
	assign leaf[580] = f[465] && !f[381] && f[297] && f[549]; // c4t404i40
	assign leaf[581] = f[465] && f[381] && !f[375] && !f[355]; // c4t404i40
	assign leaf[582] = f[465] && f[381] && !f[375] && f[355]; // c4t404i40
	assign leaf[583] = f[465] && f[381] && f[375] && !f[715]; // c4t404i40
	assign leaf[584] = f[465] && f[381] && f[375] && f[715]; // c4t404i40
	assign leaf[585] = !f[96] && !f[346] && !f[625] && !f[348]; // c4t414i41
	assign leaf[586] = !f[96] && !f[346] && !f[625] && f[348]; // c4t414i41
	assign leaf[587] = !f[96] && !f[346] && f[625] && !f[709]; // c4t414i41
	assign leaf[588] = !f[96] && !f[346] && f[625] && f[709]; // c4t414i41
	assign leaf[589] = !f[96] && f[346] && !f[340] && !f[400]; // c4t414i41
	assign leaf[590] = !f[96] && f[346] && !f[340] && f[400]; // c4t414i41
	assign leaf[591] = !f[96] && f[346] && f[340] && !f[398]; // c4t414i41
	assign leaf[592] = !f[96] && f[346] && f[340] && f[398]; // c4t414i41
	assign leaf[593] = f[96] && !f[455]; // c4t414i41
	assign leaf[594] = f[96] && f[455]; // c4t414i41
	assign leaf[595] = !f[625] && !f[491] && !f[321] && !f[411]; // c4t424i42
	assign leaf[596] = !f[625] && !f[491] && !f[321] && f[411]; // c4t424i42
	assign leaf[597] = !f[625] && !f[491] && f[321] && !f[654]; // c4t424i42
	assign leaf[598] = !f[625] && !f[491] && f[321] && f[654]; // c4t424i42
	assign leaf[599] = !f[625] && f[491] && !f[326] && !f[243]; // c4t424i42
	assign leaf[600] = !f[625] && f[491] && !f[326] && f[243]; // c4t424i42
	assign leaf[601] = !f[625] && f[491] && f[326] && !f[379]; // c4t424i42
	assign leaf[602] = !f[625] && f[491] && f[326] && f[379]; // c4t424i42
	assign leaf[603] = f[625] && !f[543] && !f[190]; // c4t424i42
	assign leaf[604] = f[625] && !f[543] && f[190] && !f[596]; // c4t424i42
	assign leaf[605] = f[625] && !f[543] && f[190] && f[596]; // c4t424i42
	assign leaf[606] = f[625] && f[543] && !f[186] && !f[268]; // c4t424i42
	assign leaf[607] = f[625] && f[543] && !f[186] && f[268]; // c4t424i42
	assign leaf[608] = f[625] && f[543] && f[186] && !f[132]; // c4t424i42
	assign leaf[609] = f[625] && f[543] && f[186] && f[132]; // c4t424i42
	assign leaf[610] = !f[398] && !f[403] && !f[181] && !f[206]; // c4t434i43
	assign leaf[611] = !f[398] && !f[403] && !f[181] && f[206]; // c4t434i43
	assign leaf[612] = !f[398] && !f[403] && f[181] && !f[184]; // c4t434i43
	assign leaf[613] = !f[398] && !f[403] && f[181] && f[184]; // c4t434i43
	assign leaf[614] = !f[398] && f[403] && !f[469] && !f[128]; // c4t434i43
	assign leaf[615] = !f[398] && f[403] && !f[469] && f[128]; // c4t434i43
	assign leaf[616] = !f[398] && f[403] && f[469] && !f[213]; // c4t434i43
	assign leaf[617] = !f[398] && f[403] && f[469] && f[213]; // c4t434i43
	assign leaf[618] = f[398] && !f[331] && !f[555] && !f[327]; // c4t434i43
	assign leaf[619] = f[398] && !f[331] && !f[555] && f[327]; // c4t434i43
	assign leaf[620] = f[398] && !f[331] && f[555] && !f[323]; // c4t434i43
	assign leaf[621] = f[398] && !f[331] && f[555] && f[323]; // c4t434i43
	assign leaf[622] = f[398] && f[331] && !f[461] && !f[382]; // c4t434i43
	assign leaf[623] = f[398] && f[331] && !f[461] && f[382]; // c4t434i43
	assign leaf[624] = f[398] && f[331] && f[461] && !f[241]; // c4t434i43
	assign leaf[625] = f[398] && f[331] && f[461] && f[241]; // c4t434i43
	assign leaf[626] = !f[102] && !f[97] && !f[714] && !f[381]; // c4t444i44
	assign leaf[627] = !f[102] && !f[97] && !f[714] && f[381]; // c4t444i44
	assign leaf[628] = !f[102] && !f[97] && f[714] && !f[237]; // c4t444i44
	assign leaf[629] = !f[102] && !f[97] && f[714] && f[237]; // c4t444i44
	assign leaf[630] = !f[102] && f[97] && !f[573]; // c4t444i44
	assign leaf[631] = !f[102] && f[97] && f[573]; // c4t444i44
	assign leaf[632] = f[102] && !f[296]; // c4t444i44
	assign leaf[633] = f[102] && f[296]; // c4t444i44
	assign leaf[634] = !f[179] && !f[635] && !f[241] && !f[158]; // c4t454i45
	assign leaf[635] = !f[179] && !f[635] && !f[241] && f[158]; // c4t454i45
	assign leaf[636] = !f[179] && !f[635] && f[241] && !f[244]; // c4t454i45
	assign leaf[637] = !f[179] && !f[635] && f[241] && f[244]; // c4t454i45
	assign leaf[638] = !f[179] && f[635] && !f[747] && !f[660]; // c4t454i45
	assign leaf[639] = !f[179] && f[635] && !f[747] && f[660]; // c4t454i45
	assign leaf[640] = !f[179] && f[635] && f[747]; // c4t454i45
	assign leaf[641] = f[179] && !f[181] && !f[204] && !f[153]; // c4t454i45
	assign leaf[642] = f[179] && !f[181] && !f[204] && f[153]; // c4t454i45
	assign leaf[643] = f[179] && !f[181] && f[204] && !f[300]; // c4t454i45
	assign leaf[644] = f[179] && !f[181] && f[204] && f[300]; // c4t454i45
	assign leaf[645] = f[179] && f[181] && !f[263] && !f[273]; // c4t454i45
	assign leaf[646] = f[179] && f[181] && !f[263] && f[273]; // c4t454i45
	assign leaf[647] = f[179] && f[181] && f[263] && !f[183]; // c4t454i45
	assign leaf[648] = f[179] && f[181] && f[263] && f[183]; // c4t454i45
	assign leaf[649] = !f[220] && !f[163] && !f[301] && !f[490]; // c4t464i46
	assign leaf[650] = !f[220] && !f[163] && !f[301] && f[490]; // c4t464i46
	assign leaf[651] = !f[220] && !f[163] && f[301] && !f[384]; // c4t464i46
	assign leaf[652] = !f[220] && !f[163] && f[301] && f[384]; // c4t464i46
	assign leaf[653] = !f[220] && f[163] && !f[187] && !f[596]; // c4t464i46
	assign leaf[654] = !f[220] && f[163] && !f[187] && f[596]; // c4t464i46
	assign leaf[655] = !f[220] && f[163] && f[187]; // c4t464i46
	assign leaf[656] = f[220] && !f[214] && !f[210] && !f[464]; // c4t464i46
	assign leaf[657] = f[220] && !f[214] && !f[210] && f[464]; // c4t464i46
	assign leaf[658] = f[220] && !f[214] && f[210] && !f[191]; // c4t464i46
	assign leaf[659] = f[220] && !f[214] && f[210] && f[191]; // c4t464i46
	assign leaf[660] = f[220] && f[214]; // c4t464i46
	assign leaf[661] = !f[744] && !f[128] && !f[404] && !f[483]; // c4t474i47
	assign leaf[662] = !f[744] && !f[128] && !f[404] && f[483]; // c4t474i47
	assign leaf[663] = !f[744] && !f[128] && f[404] && !f[496]; // c4t474i47
	assign leaf[664] = !f[744] && !f[128] && f[404] && f[496]; // c4t474i47
	assign leaf[665] = !f[744] && f[128] && !f[497] && !f[239]; // c4t474i47
	assign leaf[666] = !f[744] && f[128] && !f[497] && f[239]; // c4t474i47
	assign leaf[667] = !f[744] && f[128] && f[497] && !f[520]; // c4t474i47
	assign leaf[668] = !f[744] && f[128] && f[497] && f[520]; // c4t474i47
	assign leaf[669] = f[744] && !f[605]; // c4t474i47
	assign leaf[670] = f[744] && f[605]; // c4t474i47
	assign leaf[671] = !f[96] && !f[740] && !f[408] && !f[485]; // c4t484i48
	assign leaf[672] = !f[96] && !f[740] && !f[408] && f[485]; // c4t484i48
	assign leaf[673] = !f[96] && !f[740] && f[408] && !f[348]; // c4t484i48
	assign leaf[674] = !f[96] && !f[740] && f[408] && f[348]; // c4t484i48
	assign leaf[675] = !f[96] && f[740] && !f[234]; // c4t484i48
	assign leaf[676] = !f[96] && f[740] && f[234]; // c4t484i48
	assign leaf[677] = f[96] && !f[545]; // c4t484i48
	assign leaf[678] = f[96] && f[545]; // c4t484i48
	assign leaf[679] = !f[93] && !f[520] && !f[632] && !f[385]; // c4t494i49
	assign leaf[680] = !f[93] && !f[520] && !f[632] && f[385]; // c4t494i49
	assign leaf[681] = !f[93] && !f[520] && f[632] && !f[485]; // c4t494i49
	assign leaf[682] = !f[93] && !f[520] && f[632] && f[485]; // c4t494i49
	assign leaf[683] = !f[93] && f[520] && !f[628] && !f[236]; // c4t494i49
	assign leaf[684] = !f[93] && f[520] && !f[628] && f[236]; // c4t494i49
	assign leaf[685] = !f[93] && f[520] && f[628] && !f[241]; // c4t494i49
	assign leaf[686] = !f[93] && f[520] && f[628] && f[241]; // c4t494i49
	assign leaf[687] = f[93] && !f[456]; // c4t494i49
	assign leaf[688] = f[93] && f[456]; // c4t494i49
	assign leaf[689] = !f[286] && !f[184] && !f[240] && !f[323]; // c4t504i50
	assign leaf[690] = !f[286] && !f[184] && !f[240] && f[323]; // c4t504i50
	assign leaf[691] = !f[286] && !f[184] && f[240] && !f[238]; // c4t504i50
	assign leaf[692] = !f[286] && !f[184] && f[240] && f[238]; // c4t504i50
	assign leaf[693] = !f[286] && f[184] && !f[187] && !f[267]; // c4t504i50
	assign leaf[694] = !f[286] && f[184] && !f[187] && f[267]; // c4t504i50
	assign leaf[695] = !f[286] && f[184] && f[187] && !f[467]; // c4t504i50
	assign leaf[696] = !f[286] && f[184] && f[187] && f[467]; // c4t504i50
	assign leaf[697] = f[286] && !f[213] && !f[244] && !f[354]; // c4t504i50
	assign leaf[698] = f[286] && !f[213] && !f[244] && f[354]; // c4t504i50
	assign leaf[699] = f[286] && !f[213] && f[244] && !f[660]; // c4t504i50
	assign leaf[700] = f[286] && !f[213] && f[244] && f[660]; // c4t504i50
	assign leaf[701] = f[286] && f[213] && !f[205] && !f[687]; // c4t504i50
	assign leaf[702] = f[286] && f[213] && !f[205] && f[687]; // c4t504i50
	assign leaf[703] = f[286] && f[213] && f[205] && !f[636]; // c4t504i50
	assign leaf[704] = f[286] && f[213] && f[205] && f[636]; // c4t504i50
	assign leaf[705] = !f[397] && !f[346] && !f[348] && !f[344]; // c4t514i51
	assign leaf[706] = !f[397] && !f[346] && !f[348] && f[344]; // c4t514i51
	assign leaf[707] = !f[397] && !f[346] && f[348] && !f[490]; // c4t514i51
	assign leaf[708] = !f[397] && !f[346] && f[348] && f[490]; // c4t514i51
	assign leaf[709] = !f[397] && f[346] && !f[400] && !f[212]; // c4t514i51
	assign leaf[710] = !f[397] && f[346] && !f[400] && f[212]; // c4t514i51
	assign leaf[711] = !f[397] && f[346] && f[400] && !f[243]; // c4t514i51
	assign leaf[712] = !f[397] && f[346] && f[400] && f[243]; // c4t514i51
	assign leaf[713] = f[397] && !f[359] && !f[379] && !f[323]; // c4t514i51
	assign leaf[714] = f[397] && !f[359] && !f[379] && f[323]; // c4t514i51
	assign leaf[715] = f[397] && !f[359] && f[379] && !f[372]; // c4t514i51
	assign leaf[716] = f[397] && !f[359] && f[379] && f[372]; // c4t514i51
	assign leaf[717] = f[397] && f[359] && !f[429]; // c4t514i51
	assign leaf[718] = f[397] && f[359] && f[429]; // c4t514i51
	assign leaf[719] = !f[347] && !f[344] && !f[405] && !f[349]; // c4t524i52
	assign leaf[720] = !f[347] && !f[344] && !f[405] && f[349]; // c4t524i52
	assign leaf[721] = !f[347] && !f[344] && f[405] && !f[318]; // c4t524i52
	assign leaf[722] = !f[347] && !f[344] && f[405] && f[318]; // c4t524i52
	assign leaf[723] = !f[347] && f[344] && !f[180] && !f[264]; // c4t524i52
	assign leaf[724] = !f[347] && f[344] && !f[180] && f[264]; // c4t524i52
	assign leaf[725] = !f[347] && f[344] && f[180] && !f[661]; // c4t524i52
	assign leaf[726] = !f[347] && f[344] && f[180] && f[661]; // c4t524i52
	assign leaf[727] = f[347] && !f[341] && !f[542] && !f[240]; // c4t524i52
	assign leaf[728] = f[347] && !f[341] && !f[542] && f[240]; // c4t524i52
	assign leaf[729] = f[347] && !f[341] && f[542] && !f[526]; // c4t524i52
	assign leaf[730] = f[347] && !f[341] && f[542] && f[526]; // c4t524i52
	assign leaf[731] = f[347] && f[341] && !f[636] && !f[271]; // c4t524i52
	assign leaf[732] = f[347] && f[341] && !f[636] && f[271]; // c4t524i52
	assign leaf[733] = f[347] && f[341] && f[636]; // c4t524i52
	assign leaf[734] = !f[122] && !f[128] && !f[376] && !f[399]; // c4t534i53
	assign leaf[735] = !f[122] && !f[128] && !f[376] && f[399]; // c4t534i53
	assign leaf[736] = !f[122] && !f[128] && f[376] && !f[408]; // c4t534i53
	assign leaf[737] = !f[122] && !f[128] && f[376] && f[408]; // c4t534i53
	assign leaf[738] = !f[122] && f[128] && !f[405] && !f[598]; // c4t534i53
	assign leaf[739] = !f[122] && f[128] && !f[405] && f[598]; // c4t534i53
	assign leaf[740] = !f[122] && f[128] && f[405] && !f[267]; // c4t534i53
	assign leaf[741] = !f[122] && f[128] && f[405] && f[267]; // c4t534i53
	assign leaf[742] = f[122] && !f[546] && !f[630]; // c4t534i53
	assign leaf[743] = f[122] && !f[546] && f[630]; // c4t534i53
	assign leaf[744] = f[122] && f[546] && !f[513]; // c4t534i53
	assign leaf[745] = f[122] && f[546] && f[513]; // c4t534i53
	assign leaf[746] = !f[72] && !f[741] && !f[94] && !f[737]; // c4t544i54
	assign leaf[747] = !f[72] && !f[741] && !f[94] && f[737]; // c4t544i54
	assign leaf[748] = !f[72] && !f[741] && f[94]; // c4t544i54
	assign leaf[749] = !f[72] && f[741] && !f[264] && !f[321]; // c4t544i54
	assign leaf[750] = !f[72] && f[741] && !f[264] && f[321]; // c4t544i54
	assign leaf[751] = !f[72] && f[741] && f[264]; // c4t544i54
	assign leaf[752] = f[72]; // c4t544i54
	assign leaf[753] = !f[318] && !f[320] && !f[316] && !f[230]; // c4t554i55
	assign leaf[754] = !f[318] && !f[320] && !f[316] && f[230]; // c4t554i55
	assign leaf[755] = !f[318] && !f[320] && f[316] && !f[181]; // c4t554i55
	assign leaf[756] = !f[318] && !f[320] && f[316] && f[181]; // c4t554i55
	assign leaf[757] = !f[318] && f[320] && !f[262] && !f[347]; // c4t554i55
	assign leaf[758] = !f[318] && f[320] && !f[262] && f[347]; // c4t554i55
	assign leaf[759] = !f[318] && f[320] && f[262] && !f[633]; // c4t554i55
	assign leaf[760] = !f[318] && f[320] && f[262] && f[633]; // c4t554i55
	assign leaf[761] = f[318] && !f[321] && !f[209] && !f[265]; // c4t554i55
	assign leaf[762] = f[318] && !f[321] && !f[209] && f[265]; // c4t554i55
	assign leaf[763] = f[318] && !f[321] && f[209] && !f[212]; // c4t554i55
	assign leaf[764] = f[318] && !f[321] && f[209] && f[212]; // c4t554i55
	assign leaf[765] = f[318] && f[321] && !f[289] && !f[401]; // c4t554i55
	assign leaf[766] = f[318] && f[321] && !f[289] && f[401]; // c4t554i55
	assign leaf[767] = f[318] && f[321] && f[289] && !f[291]; // c4t554i55
	assign leaf[768] = f[318] && f[321] && f[289] && f[291]; // c4t554i55
	assign leaf[769] = !f[430] && !f[569] && !f[549] && !f[413]; // c4t564i56
	assign leaf[770] = !f[430] && !f[569] && !f[549] && f[413]; // c4t564i56
	assign leaf[771] = !f[430] && !f[569] && f[549] && !f[691]; // c4t564i56
	assign leaf[772] = !f[430] && !f[569] && f[549] && f[691]; // c4t564i56
	assign leaf[773] = !f[430] && f[569] && !f[497] && !f[680]; // c4t564i56
	assign leaf[774] = !f[430] && f[569] && !f[497] && f[680]; // c4t564i56
	assign leaf[775] = !f[430] && f[569] && f[497]; // c4t564i56
	assign leaf[776] = f[430] && !f[206] && !f[662] && !f[152]; // c4t564i56
	assign leaf[777] = f[430] && !f[206] && !f[662] && f[152]; // c4t564i56
	assign leaf[778] = f[430] && !f[206] && f[662] && !f[659]; // c4t564i56
	assign leaf[779] = f[430] && !f[206] && f[662] && f[659]; // c4t564i56
	assign leaf[780] = f[430] && f[206] && !f[237] && !f[155]; // c4t564i56
	assign leaf[781] = f[430] && f[206] && !f[237] && f[155]; // c4t564i56
	assign leaf[782] = f[430] && f[206] && f[237] && !f[272]; // c4t564i56
	assign leaf[783] = f[430] && f[206] && f[237] && f[272]; // c4t564i56
	assign leaf[784] = !f[430] && !f[300] && !f[181] && !f[265]; // c4t574i57
	assign leaf[785] = !f[430] && !f[300] && !f[181] && f[265]; // c4t574i57
	assign leaf[786] = !f[430] && !f[300] && f[181] && !f[234]; // c4t574i57
	assign leaf[787] = !f[430] && !f[300] && f[181] && f[234]; // c4t574i57
	assign leaf[788] = !f[430] && f[300] && !f[182] && !f[206]; // c4t574i57
	assign leaf[789] = !f[430] && f[300] && !f[182] && f[206]; // c4t574i57
	assign leaf[790] = !f[430] && f[300] && f[182] && !f[185]; // c4t574i57
	assign leaf[791] = !f[430] && f[300] && f[182] && f[185]; // c4t574i57
	assign leaf[792] = f[430] && !f[427] && !f[581] && !f[626]; // c4t574i57
	assign leaf[793] = f[430] && !f[427] && !f[581] && f[626]; // c4t574i57
	assign leaf[794] = f[430] && !f[427] && f[581] && !f[353]; // c4t574i57
	assign leaf[795] = f[430] && !f[427] && f[581] && f[353]; // c4t574i57
	assign leaf[796] = f[430] && f[427] && !f[513] && !f[435]; // c4t574i57
	assign leaf[797] = f[430] && f[427] && !f[513] && f[435]; // c4t574i57
	assign leaf[798] = f[430] && f[427] && f[513] && !f[497]; // c4t574i57
	assign leaf[799] = f[430] && f[427] && f[513] && f[497]; // c4t574i57
	assign leaf[800] = !f[637] && !f[286] && !f[318] && !f[320]; // c4t584i58
	assign leaf[801] = !f[637] && !f[286] && !f[318] && f[320]; // c4t584i58
	assign leaf[802] = !f[637] && !f[286] && f[318] && !f[321]; // c4t584i58
	assign leaf[803] = !f[637] && !f[286] && f[318] && f[321]; // c4t584i58
	assign leaf[804] = !f[637] && f[286] && !f[201] && !f[685]; // c4t584i58
	assign leaf[805] = !f[637] && f[286] && !f[201] && f[685]; // c4t584i58
	assign leaf[806] = !f[637] && f[286] && f[201]; // c4t584i58
	assign leaf[807] = f[637] && !f[234] && !f[151] && !f[523]; // c4t584i58
	assign leaf[808] = f[637] && !f[234] && !f[151] && f[523]; // c4t584i58
	assign leaf[809] = f[637] && !f[234] && f[151]; // c4t584i58
	assign leaf[810] = f[637] && f[234] && !f[482] && !f[462]; // c4t584i58
	assign leaf[811] = f[637] && f[234] && !f[482] && f[462]; // c4t584i58
	assign leaf[812] = f[637] && f[234] && f[482]; // c4t584i58
	assign leaf[813] = !f[743] && !f[398] && !f[347] && !f[181]; // c4t594i59
	assign leaf[814] = !f[743] && !f[398] && !f[347] && f[181]; // c4t594i59
	assign leaf[815] = !f[743] && !f[398] && f[347] && !f[313]; // c4t594i59
	assign leaf[816] = !f[743] && !f[398] && f[347] && f[313]; // c4t594i59
	assign leaf[817] = !f[743] && f[398] && !f[344] && !f[343]; // c4t594i59
	assign leaf[818] = !f[743] && f[398] && !f[344] && f[343]; // c4t594i59
	assign leaf[819] = !f[743] && f[398] && f[344] && !f[465]; // c4t594i59
	assign leaf[820] = !f[743] && f[398] && f[344] && f[465]; // c4t594i59
	assign leaf[821] = f[743] && !f[521]; // c4t594i59
	assign leaf[822] = f[743] && f[521] && !f[411]; // c4t594i59
	assign leaf[823] = f[743] && f[521] && f[411]; // c4t594i59
	assign leaf[824] = !f[179] && !f[154] && !f[404] && !f[636]; // c4t604i60
	assign leaf[825] = !f[179] && !f[154] && !f[404] && f[636]; // c4t604i60
	assign leaf[826] = !f[179] && !f[154] && f[404] && !f[434]; // c4t604i60
	assign leaf[827] = !f[179] && !f[154] && f[404] && f[434]; // c4t604i60
	assign leaf[828] = !f[179] && f[154] && !f[156] && !f[128]; // c4t604i60
	assign leaf[829] = !f[179] && f[154] && !f[156] && f[128]; // c4t604i60
	assign leaf[830] = !f[179] && f[154] && f[156] && !f[266]; // c4t604i60
	assign leaf[831] = !f[179] && f[154] && f[156] && f[266]; // c4t604i60
	assign leaf[832] = f[179] && !f[235] && !f[405] && !f[180]; // c4t604i60
	assign leaf[833] = f[179] && !f[235] && !f[405] && f[180]; // c4t604i60
	assign leaf[834] = f[179] && !f[235] && f[405] && !f[262]; // c4t604i60
	assign leaf[835] = f[179] && !f[235] && f[405] && f[262]; // c4t604i60
	assign leaf[836] = f[179] && f[235] && !f[214] && !f[181]; // c4t604i60
	assign leaf[837] = f[179] && f[235] && !f[214] && f[181]; // c4t604i60
	assign leaf[838] = f[179] && f[235] && f[214] && !f[155]; // c4t604i60
	assign leaf[839] = f[179] && f[235] && f[214] && f[155]; // c4t604i60
	assign leaf[840] = !f[519] && !f[630] && !f[686] && !f[201]; // c4t614i61
	assign leaf[841] = !f[519] && !f[630] && !f[686] && f[201]; // c4t614i61
	assign leaf[842] = !f[519] && !f[630] && f[686] && !f[660]; // c4t614i61
	assign leaf[843] = !f[519] && !f[630] && f[686] && f[660]; // c4t614i61
	assign leaf[844] = !f[519] && f[630] && !f[605] && !f[181]; // c4t614i61
	assign leaf[845] = !f[519] && f[630] && !f[605] && f[181]; // c4t614i61
	assign leaf[846] = !f[519] && f[630] && f[605] && !f[328]; // c4t614i61
	assign leaf[847] = !f[519] && f[630] && f[605] && f[328]; // c4t614i61
	assign leaf[848] = f[519] && !f[524] && !f[186] && !f[297]; // c4t614i61
	assign leaf[849] = f[519] && !f[524] && !f[186] && f[297]; // c4t614i61
	assign leaf[850] = f[519] && !f[524] && f[186] && !f[269]; // c4t614i61
	assign leaf[851] = f[519] && !f[524] && f[186] && f[269]; // c4t614i61
	assign leaf[852] = f[519] && f[524] && !f[261] && !f[387]; // c4t614i61
	assign leaf[853] = f[519] && f[524] && !f[261] && f[387]; // c4t614i61
	assign leaf[854] = f[519] && f[524] && f[261] && !f[273]; // c4t614i61
	assign leaf[855] = f[519] && f[524] && f[261] && f[273]; // c4t614i61
	assign leaf[856] = !f[318] && !f[320] && !f[316] && !f[257]; // c4t624i62
	assign leaf[857] = !f[318] && !f[320] && !f[316] && f[257]; // c4t624i62
	assign leaf[858] = !f[318] && !f[320] && f[316] && !f[264]; // c4t624i62
	assign leaf[859] = !f[318] && !f[320] && f[316] && f[264]; // c4t624i62
	assign leaf[860] = !f[318] && f[320] && !f[262] && !f[274]; // c4t624i62
	assign leaf[861] = !f[318] && f[320] && !f[262] && f[274]; // c4t624i62
	assign leaf[862] = !f[318] && f[320] && f[262] && !f[577]; // c4t624i62
	assign leaf[863] = !f[318] && f[320] && f[262] && f[577]; // c4t624i62
	assign leaf[864] = f[318] && !f[321] && !f[237] && !f[181]; // c4t624i62
	assign leaf[865] = f[318] && !f[321] && !f[237] && f[181]; // c4t624i62
	assign leaf[866] = f[318] && !f[321] && f[237] && !f[320]; // c4t624i62
	assign leaf[867] = f[318] && !f[321] && f[237] && f[320]; // c4t624i62
	assign leaf[868] = f[318] && f[321] && !f[183] && !f[289]; // c4t624i62
	assign leaf[869] = f[318] && f[321] && !f[183] && f[289]; // c4t624i62
	assign leaf[870] = f[318] && f[321] && f[183] && !f[296]; // c4t624i62
	assign leaf[871] = f[318] && f[321] && f[183] && f[296]; // c4t624i62
	assign leaf[872] = !f[381] && !f[515] && !f[321] && !f[182]; // c4t634i63
	assign leaf[873] = !f[381] && !f[515] && !f[321] && f[182]; // c4t634i63
	assign leaf[874] = !f[381] && !f[515] && f[321] && !f[662]; // c4t634i63
	assign leaf[875] = !f[381] && !f[515] && f[321] && f[662]; // c4t634i63
	assign leaf[876] = !f[381] && f[515] && !f[409] && !f[579]; // c4t634i63
	assign leaf[877] = !f[381] && f[515] && !f[409] && f[579]; // c4t634i63
	assign leaf[878] = !f[381] && f[515] && f[409] && !f[154]; // c4t634i63
	assign leaf[879] = !f[381] && f[515] && f[409] && f[154]; // c4t634i63
	assign leaf[880] = f[381] && !f[465] && !f[158] && !f[466]; // c4t634i63
	assign leaf[881] = f[381] && !f[465] && !f[158] && f[466]; // c4t634i63
	assign leaf[882] = f[381] && !f[465] && f[158] && !f[372]; // c4t634i63
	assign leaf[883] = f[381] && !f[465] && f[158] && f[372]; // c4t634i63
	assign leaf[884] = f[381] && f[465] && !f[235] && !f[316]; // c4t634i63
	assign leaf[885] = f[381] && f[465] && !f[235] && f[316]; // c4t634i63
	assign leaf[886] = f[381] && f[465] && f[235] && !f[246]; // c4t634i63
	assign leaf[887] = f[381] && f[465] && f[235] && f[246]; // c4t634i63
	assign leaf[888] = !f[128] && !f[555] && !f[348] && !f[219]; // c4t644i64
	assign leaf[889] = !f[128] && !f[555] && !f[348] && f[219]; // c4t644i64
	assign leaf[890] = !f[128] && !f[555] && f[348] && !f[716]; // c4t644i64
	assign leaf[891] = !f[128] && !f[555] && f[348] && f[716]; // c4t644i64
	assign leaf[892] = !f[128] && f[555] && !f[512] && !f[179]; // c4t644i64
	assign leaf[893] = !f[128] && f[555] && !f[512] && f[179]; // c4t644i64
	assign leaf[894] = !f[128] && f[555] && f[512]; // c4t644i64
	assign leaf[895] = f[128] && !f[405] && !f[626] && !f[126]; // c4t644i64
	assign leaf[896] = f[128] && !f[405] && !f[626] && f[126]; // c4t644i64
	assign leaf[897] = f[128] && !f[405] && f[626]; // c4t644i64
	assign leaf[898] = f[128] && f[405] && !f[129]; // c4t644i64
	assign leaf[899] = f[128] && f[405] && f[129]; // c4t644i64
	assign leaf[900] = !f[744] && !f[121] && !f[102] && !f[656]; // c4t654i65
	assign leaf[901] = !f[744] && !f[121] && !f[102] && f[656]; // c4t654i65
	assign leaf[902] = !f[744] && !f[121] && f[102] && !f[467]; // c4t654i65
	assign leaf[903] = !f[744] && !f[121] && f[102] && f[467]; // c4t654i65
	assign leaf[904] = !f[744] && f[121] && !f[484]; // c4t654i65
	assign leaf[905] = !f[744] && f[121] && f[484]; // c4t654i65
	assign leaf[906] = f[744] && !f[299]; // c4t654i65
	assign leaf[907] = f[744] && f[299]; // c4t654i65
	assign leaf[908] = !f[738] && !f[96] && !f[747] && !f[384]; // c4t664i66
	assign leaf[909] = !f[738] && !f[96] && !f[747] && f[384]; // c4t664i66
	assign leaf[910] = !f[738] && !f[96] && f[747]; // c4t664i66
	assign leaf[911] = !f[738] && f[96]; // c4t664i66
	assign leaf[912] = f[738] && !f[269]; // c4t664i66
	assign leaf[913] = f[738] && f[269]; // c4t664i66
	assign leaf[914] = !f[429] && !f[349] && !f[237] && !f[293]; // c4t674i67
	assign leaf[915] = !f[429] && !f[349] && !f[237] && f[293]; // c4t674i67
	assign leaf[916] = !f[429] && !f[349] && f[237] && !f[211]; // c4t674i67
	assign leaf[917] = !f[429] && !f[349] && f[237] && f[211]; // c4t674i67
	assign leaf[918] = !f[429] && f[349] && !f[467] && !f[454]; // c4t674i67
	assign leaf[919] = !f[429] && f[349] && !f[467] && f[454]; // c4t674i67
	assign leaf[920] = !f[429] && f[349] && f[467] && !f[184]; // c4t674i67
	assign leaf[921] = !f[429] && f[349] && f[467] && f[184]; // c4t674i67
	assign leaf[922] = f[429] && !f[205] && !f[214] && !f[210]; // c4t674i67
	assign leaf[923] = f[429] && !f[205] && !f[214] && f[210]; // c4t674i67
	assign leaf[924] = f[429] && !f[205] && f[214] && !f[272]; // c4t674i67
	assign leaf[925] = f[429] && !f[205] && f[214] && f[272]; // c4t674i67
	assign leaf[926] = f[429] && f[205] && !f[289] && !f[413]; // c4t674i67
	assign leaf[927] = f[429] && f[205] && !f[289] && f[413]; // c4t674i67
	assign leaf[928] = f[429] && f[205] && f[289] && !f[265]; // c4t674i67
	assign leaf[929] = f[429] && f[205] && f[289] && f[265]; // c4t674i67
	assign leaf[930] = !f[179] && !f[690] && !f[525] && !f[539]; // c4t684i68
	assign leaf[931] = !f[179] && !f[690] && !f[525] && f[539]; // c4t684i68
	assign leaf[932] = !f[179] && !f[690] && f[525] && !f[596]; // c4t684i68
	assign leaf[933] = !f[179] && !f[690] && f[525] && f[596]; // c4t684i68
	assign leaf[934] = !f[179] && f[690] && !f[236] && !f[239]; // c4t684i68
	assign leaf[935] = !f[179] && f[690] && !f[236] && f[239]; // c4t684i68
	assign leaf[936] = !f[179] && f[690] && f[236] && !f[181]; // c4t684i68
	assign leaf[937] = !f[179] && f[690] && f[236] && f[181]; // c4t684i68
	assign leaf[938] = f[179] && !f[263] && !f[152] && !f[181]; // c4t684i68
	assign leaf[939] = f[179] && !f[263] && !f[152] && f[181]; // c4t684i68
	assign leaf[940] = f[179] && !f[263] && f[152] && !f[483]; // c4t684i68
	assign leaf[941] = f[179] && !f[263] && f[152] && f[483]; // c4t684i68
	assign leaf[942] = f[179] && f[263] && !f[213] && !f[354]; // c4t684i68
	assign leaf[943] = f[179] && f[263] && !f[213] && f[354]; // c4t684i68
	assign leaf[944] = f[179] && f[263] && f[213] && !f[182]; // c4t684i68
	assign leaf[945] = f[179] && f[263] && f[213] && f[182]; // c4t684i68
	assign leaf[946] = !f[739] && !f[72] && !f[96] && !f[519]; // c4t694i69
	assign leaf[947] = !f[739] && !f[72] && !f[96] && f[519]; // c4t694i69
	assign leaf[948] = !f[739] && !f[72] && f[96]; // c4t694i69
	assign leaf[949] = !f[739] && f[72]; // c4t694i69
	assign leaf[950] = f[739] && !f[438]; // c4t694i69
	assign leaf[951] = f[739] && f[438]; // c4t694i69
	assign leaf[952] = !f[399] && !f[286] && !f[184] && !f[267]; // c4t704i70
	assign leaf[953] = !f[399] && !f[286] && !f[184] && f[267]; // c4t704i70
	assign leaf[954] = !f[399] && !f[286] && f[184] && !f[214]; // c4t704i70
	assign leaf[955] = !f[399] && !f[286] && f[184] && f[214]; // c4t704i70
	assign leaf[956] = !f[399] && f[286] && !f[426] && !f[211]; // c4t704i70
	assign leaf[957] = !f[399] && f[286] && !f[426] && f[211]; // c4t704i70
	assign leaf[958] = !f[399] && f[286] && f[426]; // c4t704i70
	assign leaf[959] = f[399] && !f[514] && !f[463] && !f[382]; // c4t704i70
	assign leaf[960] = f[399] && !f[514] && !f[463] && f[382]; // c4t704i70
	assign leaf[961] = f[399] && !f[514] && f[463] && !f[233]; // c4t704i70
	assign leaf[962] = f[399] && !f[514] && f[463] && f[233]; // c4t704i70
	assign leaf[963] = f[399] && f[514] && !f[467] && !f[327]; // c4t704i70
	assign leaf[964] = f[399] && f[514] && !f[467] && f[327]; // c4t704i70
	assign leaf[965] = f[399] && f[514] && f[467] && !f[382]; // c4t704i70
	assign leaf[966] = f[399] && f[514] && f[467] && f[382]; // c4t704i70
	assign leaf[967] = !f[738] && !f[741] && !f[184] && !f[240]; // c4t714i71
	assign leaf[968] = !f[738] && !f[741] && !f[184] && f[240]; // c4t714i71
	assign leaf[969] = !f[738] && !f[741] && f[184] && !f[240]; // c4t714i71
	assign leaf[970] = !f[738] && !f[741] && f[184] && f[240]; // c4t714i71
	assign leaf[971] = !f[738] && f[741] && !f[264]; // c4t714i71
	assign leaf[972] = !f[738] && f[741] && f[264]; // c4t714i71
	assign leaf[973] = f[738]; // c4t714i71
	assign leaf[974] = !f[179] && !f[153] && !f[178] && !f[263]; // c4t724i72
	assign leaf[975] = !f[179] && !f[153] && !f[178] && f[263]; // c4t724i72
	assign leaf[976] = !f[179] && !f[153] && f[178] && !f[269]; // c4t724i72
	assign leaf[977] = !f[179] && !f[153] && f[178] && f[269]; // c4t724i72
	assign leaf[978] = !f[179] && f[153] && !f[551] && !f[464]; // c4t724i72
	assign leaf[979] = !f[179] && f[153] && !f[551] && f[464]; // c4t724i72
	assign leaf[980] = !f[179] && f[153] && f[551] && !f[520]; // c4t724i72
	assign leaf[981] = !f[179] && f[153] && f[551] && f[520]; // c4t724i72
	assign leaf[982] = f[179] && !f[155] && !f[204] && !f[213]; // c4t724i72
	assign leaf[983] = f[179] && !f[155] && !f[204] && f[213]; // c4t724i72
	assign leaf[984] = f[179] && !f[155] && f[204] && !f[436]; // c4t724i72
	assign leaf[985] = f[179] && !f[155] && f[204] && f[436]; // c4t724i72
	assign leaf[986] = f[179] && f[155] && !f[540] && !f[267]; // c4t724i72
	assign leaf[987] = f[179] && f[155] && !f[540] && f[267]; // c4t724i72
	assign leaf[988] = f[179] && f[155] && f[540]; // c4t724i72
	assign leaf[989] = !f[637] && !f[444] && !f[570] && !f[624]; // c4t734i73
	assign leaf[990] = !f[637] && !f[444] && !f[570] && f[624]; // c4t734i73
	assign leaf[991] = !f[637] && !f[444] && f[570] && !f[400]; // c4t734i73
	assign leaf[992] = !f[637] && !f[444] && f[570] && f[400]; // c4t734i73
	assign leaf[993] = !f[637] && f[444] && !f[298] && !f[211]; // c4t734i73
	assign leaf[994] = !f[637] && f[444] && !f[298] && f[211]; // c4t734i73
	assign leaf[995] = !f[637] && f[444] && f[298] && !f[454]; // c4t734i73
	assign leaf[996] = !f[637] && f[444] && f[298] && f[454]; // c4t734i73
	assign leaf[997] = f[637] && !f[234] && !f[522]; // c4t734i73
	assign leaf[998] = f[637] && !f[234] && f[522] && !f[399]; // c4t734i73
	assign leaf[999] = f[637] && !f[234] && f[522] && f[399]; // c4t734i73
	assign leaf[1000] = f[637] && f[234] && !f[453] && !f[210]; // c4t734i73
	assign leaf[1001] = f[637] && f[234] && !f[453] && f[210]; // c4t734i73
	assign leaf[1002] = f[637] && f[234] && f[453]; // c4t734i73
	assign leaf[1003] = !f[601] && !f[657] && !f[441] && !f[459]; // c4t744i74
	assign leaf[1004] = !f[601] && !f[657] && !f[441] && f[459]; // c4t744i74
	assign leaf[1005] = !f[601] && !f[657] && f[441] && !f[217]; // c4t744i74
	assign leaf[1006] = !f[601] && !f[657] && f[441] && f[217]; // c4t744i74
	assign leaf[1007] = !f[601] && f[657] && !f[437] && !f[267]; // c4t744i74
	assign leaf[1008] = !f[601] && f[657] && !f[437] && f[267]; // c4t744i74
	assign leaf[1009] = !f[601] && f[657] && f[437] && !f[547]; // c4t744i74
	assign leaf[1010] = !f[601] && f[657] && f[437] && f[547]; // c4t744i74
	assign leaf[1011] = f[601] && !f[518] && !f[399]; // c4t744i74
	assign leaf[1012] = f[601] && !f[518] && f[399] && !f[240]; // c4t744i74
	assign leaf[1013] = f[601] && !f[518] && f[399] && f[240]; // c4t744i74
	assign leaf[1014] = f[601] && f[518] && !f[239] && !f[322]; // c4t744i74
	assign leaf[1015] = f[601] && f[518] && !f[239] && f[322]; // c4t744i74
	assign leaf[1016] = f[601] && f[518] && f[239] && !f[468]; // c4t744i74
	assign leaf[1017] = f[601] && f[518] && f[239] && f[468]; // c4t744i74
	assign leaf[1018] = !f[737] && !f[303] && !f[398] && !f[347]; // c4t754i75
	assign leaf[1019] = !f[737] && !f[303] && !f[398] && f[347]; // c4t754i75
	assign leaf[1020] = !f[737] && !f[303] && f[398] && !f[294]; // c4t754i75
	assign leaf[1021] = !f[737] && !f[303] && f[398] && f[294]; // c4t754i75
	assign leaf[1022] = !f[737] && f[303] && !f[453] && !f[324]; // c4t754i75
	assign leaf[1023] = !f[737] && f[303] && !f[453] && f[324]; // c4t754i75
	assign leaf[1024] = !f[737] && f[303] && f[453]; // c4t754i75
	assign leaf[1025] = f[737]; // c4t754i75
	assign leaf[1026] = !f[746] && !f[376] && !f[321] && !f[182]; // c4t764i76
	assign leaf[1027] = !f[746] && !f[376] && !f[321] && f[182]; // c4t764i76
	assign leaf[1028] = !f[746] && !f[376] && f[321] && !f[238]; // c4t764i76
	assign leaf[1029] = !f[746] && !f[376] && f[321] && f[238]; // c4t764i76
	assign leaf[1030] = !f[746] && f[376] && !f[435] && !f[296]; // c4t764i76
	assign leaf[1031] = !f[746] && f[376] && !f[435] && f[296]; // c4t764i76
	assign leaf[1032] = !f[746] && f[376] && f[435] && !f[155]; // c4t764i76
	assign leaf[1033] = !f[746] && f[376] && f[435] && f[155]; // c4t764i76
	assign leaf[1034] = f[746]; // c4t764i76
	assign leaf[1035] = !f[465] && !f[238] && !f[213] && !f[215]; // c4t774i77
	assign leaf[1036] = !f[465] && !f[238] && !f[213] && f[215]; // c4t774i77
	assign leaf[1037] = !f[465] && !f[238] && f[213] && !f[182]; // c4t774i77
	assign leaf[1038] = !f[465] && !f[238] && f[213] && f[182]; // c4t774i77
	assign leaf[1039] = !f[465] && f[238] && !f[240] && !f[186]; // c4t774i77
	assign leaf[1040] = !f[465] && f[238] && !f[240] && f[186]; // c4t774i77
	assign leaf[1041] = !f[465] && f[238] && f[240] && !f[242]; // c4t774i77
	assign leaf[1042] = !f[465] && f[238] && f[240] && f[242]; // c4t774i77
	assign leaf[1043] = f[465] && !f[340] && !f[242] && !f[328]; // c4t774i77
	assign leaf[1044] = f[465] && !f[340] && !f[242] && f[328]; // c4t774i77
	assign leaf[1045] = f[465] && !f[340] && f[242] && !f[328]; // c4t774i77
	assign leaf[1046] = f[465] && !f[340] && f[242] && f[328]; // c4t774i77
	assign leaf[1047] = f[465] && f[340] && !f[240] && !f[352]; // c4t774i77
	assign leaf[1048] = f[465] && f[340] && !f[240] && f[352]; // c4t774i77
	assign leaf[1049] = f[465] && f[340] && f[240]; // c4t774i77
	assign leaf[1050] = !f[102] && !f[430] && !f[379] && !f[580]; // c4t784i78
	assign leaf[1051] = !f[102] && !f[430] && !f[379] && f[580]; // c4t784i78
	assign leaf[1052] = !f[102] && !f[430] && f[379] && !f[459]; // c4t784i78
	assign leaf[1053] = !f[102] && !f[430] && f[379] && f[459]; // c4t784i78
	assign leaf[1054] = !f[102] && f[430] && !f[709] && !f[579]; // c4t784i78
	assign leaf[1055] = !f[102] && f[430] && !f[709] && f[579]; // c4t784i78
	assign leaf[1056] = !f[102] && f[430] && f[709] && !f[570]; // c4t784i78
	assign leaf[1057] = !f[102] && f[430] && f[709] && f[570]; // c4t784i78
	assign leaf[1058] = f[102] && !f[185]; // c4t784i78
	assign leaf[1059] = f[102] && f[185]; // c4t784i78
	assign leaf[1060] = !f[685] && !f[320] && !f[289] && !f[287]; // c4t794i79
	assign leaf[1061] = !f[685] && !f[320] && !f[289] && f[287]; // c4t794i79
	assign leaf[1062] = !f[685] && !f[320] && f[289] && !f[180]; // c4t794i79
	assign leaf[1063] = !f[685] && !f[320] && f[289] && f[180]; // c4t794i79
	assign leaf[1064] = !f[685] && f[320] && !f[237] && !f[211]; // c4t794i79
	assign leaf[1065] = !f[685] && f[320] && !f[237] && f[211]; // c4t794i79
	assign leaf[1066] = !f[685] && f[320] && f[237] && !f[289]; // c4t794i79
	assign leaf[1067] = !f[685] && f[320] && f[237] && f[289]; // c4t794i79
	assign leaf[1068] = f[685] && !f[239] && !f[184] && !f[322]; // c4t794i79
	assign leaf[1069] = f[685] && !f[239] && !f[184] && f[322]; // c4t794i79
	assign leaf[1070] = f[685] && !f[239] && f[184] && !f[183]; // c4t794i79
	assign leaf[1071] = f[685] && !f[239] && f[184] && f[183]; // c4t794i79
	assign leaf[1072] = f[685] && f[239] && !f[322] && !f[433]; // c4t794i79
	assign leaf[1073] = f[685] && f[239] && !f[322] && f[433]; // c4t794i79
	assign leaf[1074] = f[685] && f[239] && f[322] && !f[460]; // c4t794i79
	assign leaf[1075] = f[685] && f[239] && f[322] && f[460]; // c4t794i79
	assign leaf[1076] = !f[385] && !f[320] && !f[237] && !f[181]; // c4t804i80
	assign leaf[1077] = !f[385] && !f[320] && !f[237] && f[181]; // c4t804i80
	assign leaf[1078] = !f[385] && !f[320] && f[237] && !f[154]; // c4t804i80
	assign leaf[1079] = !f[385] && !f[320] && f[237] && f[154]; // c4t804i80
	assign leaf[1080] = !f[385] && f[320] && !f[152] && !f[162]; // c4t804i80
	assign leaf[1081] = !f[385] && f[320] && !f[152] && f[162]; // c4t804i80
	assign leaf[1082] = !f[385] && f[320] && f[152] && !f[600]; // c4t804i80
	assign leaf[1083] = !f[385] && f[320] && f[152] && f[600]; // c4t804i80
	assign leaf[1084] = f[385] && !f[522] && !f[539] && !f[435]; // c4t804i80
	assign leaf[1085] = f[385] && !f[522] && !f[539] && f[435]; // c4t804i80
	assign leaf[1086] = f[385] && !f[522] && f[539] && !f[345]; // c4t804i80
	assign leaf[1087] = f[385] && !f[522] && f[539] && f[345]; // c4t804i80
	assign leaf[1088] = f[385] && f[522] && !f[353] && !f[464]; // c4t804i80
	assign leaf[1089] = f[385] && f[522] && !f[353] && f[464]; // c4t804i80
	assign leaf[1090] = f[385] && f[522] && f[353] && !f[518]; // c4t804i80
	assign leaf[1091] = f[385] && f[522] && f[353] && f[518]; // c4t804i80
	assign leaf[1092] = !f[121] && !f[186] && !f[188] && !f[269]; // c4t814i81
	assign leaf[1093] = !f[121] && !f[186] && !f[188] && f[269]; // c4t814i81
	assign leaf[1094] = !f[121] && !f[186] && f[188] && !f[601]; // c4t814i81
	assign leaf[1095] = !f[121] && !f[186] && f[188] && f[601]; // c4t814i81
	assign leaf[1096] = !f[121] && f[186] && !f[269] && !f[295]; // c4t814i81
	assign leaf[1097] = !f[121] && f[186] && !f[269] && f[295]; // c4t814i81
	assign leaf[1098] = !f[121] && f[186] && f[269] && !f[469]; // c4t814i81
	assign leaf[1099] = !f[121] && f[186] && f[269] && f[469]; // c4t814i81
	assign leaf[1100] = f[121] && !f[574]; // c4t814i81
	assign leaf[1101] = f[121] && f[574]; // c4t814i81
	assign leaf[1102] = !f[738] && !f[72] && !f[94] && !f[383]; // c4t824i82
	assign leaf[1103] = !f[738] && !f[72] && !f[94] && f[383]; // c4t824i82
	assign leaf[1104] = !f[738] && !f[72] && f[94]; // c4t824i82
	assign leaf[1105] = !f[738] && f[72]; // c4t824i82
	assign leaf[1106] = f[738]; // c4t824i82
	assign leaf[1107] = !f[384] && !f[494] && !f[435] && !f[294]; // c4t834i83
	assign leaf[1108] = !f[384] && !f[494] && !f[435] && f[294]; // c4t834i83
	assign leaf[1109] = !f[384] && !f[494] && f[435] && !f[326]; // c4t834i83
	assign leaf[1110] = !f[384] && !f[494] && f[435] && f[326]; // c4t834i83
	assign leaf[1111] = !f[384] && f[494] && !f[206] && !f[518]; // c4t834i83
	assign leaf[1112] = !f[384] && f[494] && !f[206] && f[518]; // c4t834i83
	assign leaf[1113] = !f[384] && f[494] && f[206] && !f[210]; // c4t834i83
	assign leaf[1114] = !f[384] && f[494] && f[206] && f[210]; // c4t834i83
	assign leaf[1115] = f[384] && !f[439] && !f[486] && !f[351]; // c4t834i83
	assign leaf[1116] = f[384] && !f[439] && !f[486] && f[351]; // c4t834i83
	assign leaf[1117] = f[384] && !f[439] && f[486] && !f[210]; // c4t834i83
	assign leaf[1118] = f[384] && !f[439] && f[486] && f[210]; // c4t834i83
	assign leaf[1119] = f[384] && f[439] && !f[353] && !f[214]; // c4t834i83
	assign leaf[1120] = f[384] && f[439] && !f[353] && f[214]; // c4t834i83
	assign leaf[1121] = f[384] && f[439] && f[353] && !f[271]; // c4t834i83
	assign leaf[1122] = f[384] && f[439] && f[353] && f[271]; // c4t834i83
	assign leaf[1123] = !f[275] && !f[123] && !f[238] && !f[240]; // c4t844i84
	assign leaf[1124] = !f[275] && !f[123] && !f[238] && f[240]; // c4t844i84
	assign leaf[1125] = !f[275] && !f[123] && f[238] && !f[154]; // c4t844i84
	assign leaf[1126] = !f[275] && !f[123] && f[238] && f[154]; // c4t844i84
	assign leaf[1127] = !f[275] && f[123] && !f[484]; // c4t844i84
	assign leaf[1128] = !f[275] && f[123] && f[484]; // c4t844i84
	assign leaf[1129] = f[275] && !f[453] && !f[385] && !f[237]; // c4t844i84
	assign leaf[1130] = f[275] && !f[453] && !f[385] && f[237]; // c4t844i84
	assign leaf[1131] = f[275] && !f[453] && f[385] && !f[245]; // c4t844i84
	assign leaf[1132] = f[275] && !f[453] && f[385] && f[245]; // c4t844i84
	assign leaf[1133] = f[275] && f[453]; // c4t844i84
	assign leaf[1134] = !f[663] && !f[606] && !f[579] && !f[513]; // c4t854i85
	assign leaf[1135] = !f[663] && !f[606] && !f[579] && f[513]; // c4t854i85
	assign leaf[1136] = !f[663] && !f[606] && f[579] && !f[213]; // c4t854i85
	assign leaf[1137] = !f[663] && !f[606] && f[579] && f[213]; // c4t854i85
	assign leaf[1138] = !f[663] && f[606] && !f[549]; // c4t854i85
	assign leaf[1139] = !f[663] && f[606] && f[549] && !f[349]; // c4t854i85
	assign leaf[1140] = !f[663] && f[606] && f[549] && f[349]; // c4t854i85
	assign leaf[1141] = f[663] && !f[462] && !f[267] && !f[578]; // c4t854i85
	assign leaf[1142] = f[663] && !f[462] && !f[267] && f[578]; // c4t854i85
	assign leaf[1143] = f[663] && !f[462] && f[267] && !f[464]; // c4t854i85
	assign leaf[1144] = f[663] && !f[462] && f[267] && f[464]; // c4t854i85
	assign leaf[1145] = f[663] && f[462] && !f[206] && !f[290]; // c4t854i85
	assign leaf[1146] = f[663] && f[462] && !f[206] && f[290]; // c4t854i85
	assign leaf[1147] = f[663] && f[462] && f[206] && !f[232]; // c4t854i85
	assign leaf[1148] = f[663] && f[462] && f[206] && f[232]; // c4t854i85
	assign leaf[1149] = !f[184] && !f[182] && !f[294] && !f[239]; // c4t864i86
	assign leaf[1150] = !f[184] && !f[182] && !f[294] && f[239]; // c4t864i86
	assign leaf[1151] = !f[184] && !f[182] && f[294] && !f[291]; // c4t864i86
	assign leaf[1152] = !f[184] && !f[182] && f[294] && f[291]; // c4t864i86
	assign leaf[1153] = !f[184] && f[182] && !f[206] && !f[294]; // c4t864i86
	assign leaf[1154] = !f[184] && f[182] && !f[206] && f[294]; // c4t864i86
	assign leaf[1155] = !f[184] && f[182] && f[206] && !f[291]; // c4t864i86
	assign leaf[1156] = !f[184] && f[182] && f[206] && f[291]; // c4t864i86
	assign leaf[1157] = f[184] && !f[215] && !f[239] && !f[268]; // c4t864i86
	assign leaf[1158] = f[184] && !f[215] && !f[239] && f[268]; // c4t864i86
	assign leaf[1159] = f[184] && !f[215] && f[239] && !f[159]; // c4t864i86
	assign leaf[1160] = f[184] && !f[215] && f[239] && f[159]; // c4t864i86
	assign leaf[1161] = f[184] && f[215] && !f[581] && !f[441]; // c4t864i86
	assign leaf[1162] = f[184] && f[215] && !f[581] && f[441]; // c4t864i86
	assign leaf[1163] = f[184] && f[215] && f[581]; // c4t864i86
	assign leaf[1164] = !f[746] && !f[429] && !f[349] && !f[188]; // c4t874i87
	assign leaf[1165] = !f[746] && !f[429] && !f[349] && f[188]; // c4t874i87
	assign leaf[1166] = !f[746] && !f[429] && f[349] && !f[466]; // c4t874i87
	assign leaf[1167] = !f[746] && !f[429] && f[349] && f[466]; // c4t874i87
	assign leaf[1168] = !f[746] && f[429] && !f[397] && !f[374]; // c4t874i87
	assign leaf[1169] = !f[746] && f[429] && !f[397] && f[374]; // c4t874i87
	assign leaf[1170] = !f[746] && f[429] && f[397] && !f[382]; // c4t874i87
	assign leaf[1171] = !f[746] && f[429] && f[397] && f[382]; // c4t874i87
	assign leaf[1172] = f[746]; // c4t874i87
	assign leaf[1173] = !f[465] && !f[424] && !f[380] && !f[439]; // c4t884i88
	assign leaf[1174] = !f[465] && !f[424] && !f[380] && f[439]; // c4t884i88
	assign leaf[1175] = !f[465] && !f[424] && f[380] && !f[466]; // c4t884i88
	assign leaf[1176] = !f[465] && !f[424] && f[380] && f[466]; // c4t884i88
	assign leaf[1177] = !f[465] && f[424]; // c4t884i88
	assign leaf[1178] = f[465] && !f[431] && !f[467] && !f[316]; // c4t884i88
	assign leaf[1179] = f[465] && !f[431] && !f[467] && f[316]; // c4t884i88
	assign leaf[1180] = f[465] && !f[431] && f[467] && !f[427]; // c4t884i88
	assign leaf[1181] = f[465] && !f[431] && f[467] && f[427]; // c4t884i88
	assign leaf[1182] = f[465] && f[431] && !f[216] && !f[286]; // c4t884i88
	assign leaf[1183] = f[465] && f[431] && !f[216] && f[286]; // c4t884i88
	assign leaf[1184] = f[465] && f[431] && f[216] && !f[184]; // c4t884i88
	assign leaf[1185] = f[465] && f[431] && f[216] && f[184]; // c4t884i88
	assign leaf[1186] = !f[303] && !f[386] && !f[234] && !f[684]; // c4t894i89
	assign leaf[1187] = !f[303] && !f[386] && !f[234] && f[684]; // c4t894i89
	assign leaf[1188] = !f[303] && !f[386] && f[234] && !f[237]; // c4t894i89
	assign leaf[1189] = !f[303] && !f[386] && f[234] && f[237]; // c4t894i89
	assign leaf[1190] = !f[303] && f[386] && !f[441] && !f[240]; // c4t894i89
	assign leaf[1191] = !f[303] && f[386] && !f[441] && f[240]; // c4t894i89
	assign leaf[1192] = !f[303] && f[386] && f[441] && !f[581]; // c4t894i89
	assign leaf[1193] = !f[303] && f[386] && f[441] && f[581]; // c4t894i89
	assign leaf[1194] = f[303] && !f[324] && !f[216] && !f[399]; // c4t894i89
	assign leaf[1195] = f[303] && !f[324] && !f[216] && f[399]; // c4t894i89
	assign leaf[1196] = f[303] && !f[324] && f[216]; // c4t894i89
	assign leaf[1197] = f[303] && f[324]; // c4t894i89
	assign leaf[1198] = !f[389] && !f[128] && !f[555] && !f[370]; // c4t904i90
	assign leaf[1199] = !f[389] && !f[128] && !f[555] && f[370]; // c4t904i90
	assign leaf[1200] = !f[389] && !f[128] && f[555] && !f[466]; // c4t904i90
	assign leaf[1201] = !f[389] && !f[128] && f[555] && f[466]; // c4t904i90
	assign leaf[1202] = !f[389] && f[128] && !f[497] && !f[376]; // c4t904i90
	assign leaf[1203] = !f[389] && f[128] && !f[497] && f[376]; // c4t904i90
	assign leaf[1204] = !f[389] && f[128] && f[497] && !f[293]; // c4t904i90
	assign leaf[1205] = !f[389] && f[128] && f[497] && f[293]; // c4t904i90
	assign leaf[1206] = f[389]; // c4t904i90
	assign leaf[1207] = !f[746] && !f[400] && !f[490] && !f[628]; // c4t914i91
	assign leaf[1208] = !f[746] && !f[400] && !f[490] && f[628]; // c4t914i91
	assign leaf[1209] = !f[746] && !f[400] && f[490] && !f[376]; // c4t914i91
	assign leaf[1210] = !f[746] && !f[400] && f[490] && f[376]; // c4t914i91
	assign leaf[1211] = !f[746] && f[400] && !f[547] && !f[658]; // c4t914i91
	assign leaf[1212] = !f[746] && f[400] && !f[547] && f[658]; // c4t914i91
	assign leaf[1213] = !f[746] && f[400] && f[547] && !f[549]; // c4t914i91
	assign leaf[1214] = !f[746] && f[400] && f[547] && f[549]; // c4t914i91
	assign leaf[1215] = f[746]; // c4t914i91
	assign leaf[1216] = !f[494] && !f[435] && !f[520] && !f[408]; // c4t924i92
	assign leaf[1217] = !f[494] && !f[435] && !f[520] && f[408]; // c4t924i92
	assign leaf[1218] = !f[494] && !f[435] && f[520] && !f[295]; // c4t924i92
	assign leaf[1219] = !f[494] && !f[435] && f[520] && f[295]; // c4t924i92
	assign leaf[1220] = !f[494] && f[435] && !f[238] && !f[264]; // c4t924i92
	assign leaf[1221] = !f[494] && f[435] && !f[238] && f[264]; // c4t924i92
	assign leaf[1222] = !f[494] && f[435] && f[238] && !f[294]; // c4t924i92
	assign leaf[1223] = !f[494] && f[435] && f[238] && f[294]; // c4t924i92
	assign leaf[1224] = f[494] && !f[434] && !f[350] && !f[600]; // c4t924i92
	assign leaf[1225] = f[494] && !f[434] && !f[350] && f[600]; // c4t924i92
	assign leaf[1226] = f[494] && !f[434] && f[350] && !f[635]; // c4t924i92
	assign leaf[1227] = f[494] && !f[434] && f[350] && f[635]; // c4t924i92
	assign leaf[1228] = f[494] && f[434] && !f[510] && !f[454]; // c4t924i92
	assign leaf[1229] = f[494] && f[434] && !f[510] && f[454]; // c4t924i92
	assign leaf[1230] = f[494] && f[434] && f[510] && !f[498]; // c4t924i92
	assign leaf[1231] = f[494] && f[434] && f[510] && f[498]; // c4t924i92
	assign leaf[1232] = !f[237] && !f[261] && !f[239] && !f[236]; // c4t934i93
	assign leaf[1233] = !f[237] && !f[261] && !f[239] && f[236]; // c4t934i93
	assign leaf[1234] = !f[237] && !f[261] && f[239] && !f[215]; // c4t934i93
	assign leaf[1235] = !f[237] && !f[261] && f[239] && f[215]; // c4t934i93
	assign leaf[1236] = !f[237] && f[261] && !f[181] && !f[265]; // c4t934i93
	assign leaf[1237] = !f[237] && f[261] && !f[181] && f[265]; // c4t934i93
	assign leaf[1238] = !f[237] && f[261] && f[181] && !f[629]; // c4t934i93
	assign leaf[1239] = !f[237] && f[261] && f[181] && f[629]; // c4t934i93
	assign leaf[1240] = f[237] && !f[261] && !f[185] && !f[271]; // c4t934i93
	assign leaf[1241] = f[237] && !f[261] && !f[185] && f[271]; // c4t934i93
	assign leaf[1242] = f[237] && !f[261] && f[185] && !f[215]; // c4t934i93
	assign leaf[1243] = f[237] && !f[261] && f[185] && f[215]; // c4t934i93
	assign leaf[1244] = f[237] && f[261] && !f[272] && !f[663]; // c4t934i93
	assign leaf[1245] = f[237] && f[261] && !f[272] && f[663]; // c4t934i93
	assign leaf[1246] = f[237] && f[261] && f[272] && !f[241]; // c4t934i93
	assign leaf[1247] = f[237] && f[261] && f[272] && f[241]; // c4t934i93
	assign leaf[1248] = !f[234] && !f[178] && !f[232] && !f[180]; // c4t944i94
	assign leaf[1249] = !f[234] && !f[178] && !f[232] && f[180]; // c4t944i94
	assign leaf[1250] = !f[234] && !f[178] && f[232] && !f[544]; // c4t944i94
	assign leaf[1251] = !f[234] && !f[178] && f[232] && f[544]; // c4t944i94
	assign leaf[1252] = !f[234] && f[178] && !f[179]; // c4t944i94
	assign leaf[1253] = !f[234] && f[178] && f[179] && !f[352]; // c4t944i94
	assign leaf[1254] = !f[234] && f[178] && f[179] && f[352]; // c4t944i94
	assign leaf[1255] = f[234] && !f[290] && !f[273] && !f[150]; // c4t944i94
	assign leaf[1256] = f[234] && !f[290] && !f[273] && f[150]; // c4t944i94
	assign leaf[1257] = f[234] && !f[290] && f[273]; // c4t944i94
	assign leaf[1258] = f[234] && f[290] && !f[209] && !f[239]; // c4t944i94
	assign leaf[1259] = f[234] && f[290] && !f[209] && f[239]; // c4t944i94
	assign leaf[1260] = f[234] && f[290] && f[209] && !f[239]; // c4t944i94
	assign leaf[1261] = f[234] && f[290] && f[209] && f[239]; // c4t944i94
	assign leaf[1262] = !f[741] && !f[97] && !f[381] && !f[379]; // c4t954i95
	assign leaf[1263] = !f[741] && !f[97] && !f[381] && f[379]; // c4t954i95
	assign leaf[1264] = !f[741] && !f[97] && f[381] && !f[373]; // c4t954i95
	assign leaf[1265] = !f[741] && !f[97] && f[381] && f[373]; // c4t954i95
	assign leaf[1266] = !f[741] && f[97]; // c4t954i95
	assign leaf[1267] = f[741] && !f[462]; // c4t954i95
	assign leaf[1268] = f[741] && f[462]; // c4t954i95
	assign leaf[1269] = !f[400] && !f[349] && !f[211] && !f[294]; // c4t964i96
	assign leaf[1270] = !f[400] && !f[349] && !f[211] && f[294]; // c4t964i96
	assign leaf[1271] = !f[400] && !f[349] && f[211] && !f[237]; // c4t964i96
	assign leaf[1272] = !f[400] && !f[349] && f[211] && f[237]; // c4t964i96
	assign leaf[1273] = !f[400] && f[349] && !f[179] && !f[319]; // c4t964i96
	assign leaf[1274] = !f[400] && f[349] && !f[179] && f[319]; // c4t964i96
	assign leaf[1275] = !f[400] && f[349] && f[179] && !f[206]; // c4t964i96
	assign leaf[1276] = !f[400] && f[349] && f[179] && f[206]; // c4t964i96
	assign leaf[1277] = f[400] && !f[457] && !f[628] && !f[213]; // c4t964i96
	assign leaf[1278] = f[400] && !f[457] && !f[628] && f[213]; // c4t964i96
	assign leaf[1279] = f[400] && !f[457] && f[628] && !f[517]; // c4t964i96
	assign leaf[1280] = f[400] && !f[457] && f[628] && f[517]; // c4t964i96
	assign leaf[1281] = f[400] && f[457] && !f[439] && !f[437]; // c4t964i96
	assign leaf[1282] = f[400] && f[457] && !f[439] && f[437]; // c4t964i96
	assign leaf[1283] = f[400] && f[457] && f[439] && !f[520]; // c4t964i96
	assign leaf[1284] = f[400] && f[457] && f[439] && f[520]; // c4t964i96
	assign leaf[1285] = !f[708] && !f[267] && !f[184] && !f[215]; // c4t974i97
	assign leaf[1286] = !f[708] && !f[267] && !f[184] && f[215]; // c4t974i97
	assign leaf[1287] = !f[708] && !f[267] && f[184] && !f[268]; // c4t974i97
	assign leaf[1288] = !f[708] && !f[267] && f[184] && f[268]; // c4t974i97
	assign leaf[1289] = !f[708] && f[267] && !f[242] && !f[236]; // c4t974i97
	assign leaf[1290] = !f[708] && f[267] && !f[242] && f[236]; // c4t974i97
	assign leaf[1291] = !f[708] && f[267] && f[242] && !f[497]; // c4t974i97
	assign leaf[1292] = !f[708] && f[267] && f[242] && f[497]; // c4t974i97
	assign leaf[1293] = f[708] && !f[241]; // c4t974i97
	assign leaf[1294] = f[708] && f[241]; // c4t974i97
	assign leaf[1295] = !f[637] && !f[409] && !f[681] && !f[398]; // c4t984i98
	assign leaf[1296] = !f[637] && !f[409] && !f[681] && f[398]; // c4t984i98
	assign leaf[1297] = !f[637] && !f[409] && f[681]; // c4t984i98
	assign leaf[1298] = !f[637] && f[409] && !f[348] && !f[401]; // c4t984i98
	assign leaf[1299] = !f[637] && f[409] && !f[348] && f[401]; // c4t984i98
	assign leaf[1300] = !f[637] && f[409] && f[348] && !f[296]; // c4t984i98
	assign leaf[1301] = !f[637] && f[409] && f[348] && f[296]; // c4t984i98
	assign leaf[1302] = f[637] && !f[205] && !f[523]; // c4t984i98
	assign leaf[1303] = f[637] && !f[205] && f[523] && !f[435]; // c4t984i98
	assign leaf[1304] = f[637] && !f[205] && f[523] && f[435]; // c4t984i98
	assign leaf[1305] = f[637] && f[205] && !f[180]; // c4t984i98
	assign leaf[1306] = f[637] && f[205] && f[180]; // c4t984i98
	assign leaf[1307] = !f[102] && !f[432] && !f[523] && !f[233]; // c4t994i99
	assign leaf[1308] = !f[102] && !f[432] && !f[523] && f[233]; // c4t994i99
	assign leaf[1309] = !f[102] && !f[432] && f[523] && !f[635]; // c4t994i99
	assign leaf[1310] = !f[102] && !f[432] && f[523] && f[635]; // c4t994i99
	assign leaf[1311] = !f[102] && f[432] && !f[511] && !f[232]; // c4t994i99
	assign leaf[1312] = !f[102] && f[432] && !f[511] && f[232]; // c4t994i99
	assign leaf[1313] = !f[102] && f[432] && f[511] && !f[515]; // c4t994i99
	assign leaf[1314] = !f[102] && f[432] && f[511] && f[515]; // c4t994i99
	assign leaf[1315] = f[102]; // c4t994i99
endmodule

module decision_tree_leaves_5(input logic [0:783] f, output logic [0:1401] leaf);
	assign leaf[0] = !f[220] && !f[163] && !f[276] && !f[347]; // c5t5i0
	assign leaf[1] = !f[220] && !f[163] && !f[276] && f[347]; // c5t5i0
	assign leaf[2] = !f[220] && !f[163] && f[276] && !f[330]; // c5t5i0
	assign leaf[3] = !f[220] && !f[163] && f[276] && f[330]; // c5t5i0
	assign leaf[4] = !f[220] && f[163] && !f[272] && !f[302]; // c5t5i0
	assign leaf[5] = !f[220] && f[163] && !f[272] && f[302]; // c5t5i0
	assign leaf[6] = !f[220] && f[163] && f[272] && !f[299]; // c5t5i0
	assign leaf[7] = !f[220] && f[163] && f[272] && f[299]; // c5t5i0
	assign leaf[8] = f[220] && !f[328] && !f[358] && !f[326]; // c5t5i0
	assign leaf[9] = f[220] && !f[328] && !f[358] && f[326]; // c5t5i0
	assign leaf[10] = f[220] && !f[328] && f[358]; // c5t5i0
	assign leaf[11] = f[220] && f[328] && !f[355] && !f[276]; // c5t5i0
	assign leaf[12] = f[220] && f[328] && !f[355] && f[276]; // c5t5i0
	assign leaf[13] = f[220] && f[328] && f[355] && !f[382]; // c5t5i0
	assign leaf[14] = f[220] && f[328] && f[355] && f[382]; // c5t5i0
	assign leaf[15] = !f[347] && !f[248] && !f[192] && !f[375]; // c5t15i1
	assign leaf[16] = !f[347] && !f[248] && !f[192] && f[375]; // c5t15i1
	assign leaf[17] = !f[347] && !f[248] && f[192] && !f[300]; // c5t15i1
	assign leaf[18] = !f[347] && !f[248] && f[192] && f[300]; // c5t15i1
	assign leaf[19] = !f[347] && f[248] && !f[355] && !f[359]; // c5t15i1
	assign leaf[20] = !f[347] && f[248] && !f[355] && f[359]; // c5t15i1
	assign leaf[21] = !f[347] && f[248] && f[355]; // c5t15i1
	assign leaf[22] = f[347] && !f[326] && !f[515] && !f[329]; // c5t15i1
	assign leaf[23] = f[347] && !f[326] && !f[515] && f[329]; // c5t15i1
	assign leaf[24] = f[347] && !f[326] && f[515] && !f[247]; // c5t15i1
	assign leaf[25] = f[347] && !f[326] && f[515] && f[247]; // c5t15i1
	assign leaf[26] = f[347] && f[326] && !f[408] && !f[270]; // c5t15i1
	assign leaf[27] = f[347] && f[326] && !f[408] && f[270]; // c5t15i1
	assign leaf[28] = f[347] && f[326] && f[408] && !f[304]; // c5t15i1
	assign leaf[29] = f[347] && f[326] && f[408] && f[304]; // c5t15i1
	assign leaf[30] = !f[326] && !f[296] && !f[356] && !f[655]; // c5t25i2
	assign leaf[31] = !f[326] && !f[296] && !f[356] && f[655]; // c5t25i2
	assign leaf[32] = !f[326] && !f[296] && f[356] && !f[351]; // c5t25i2
	assign leaf[33] = !f[326] && !f[296] && f[356] && f[351]; // c5t25i2
	assign leaf[34] = !f[326] && f[296] && !f[246] && !f[275]; // c5t25i2
	assign leaf[35] = !f[326] && f[296] && !f[246] && f[275]; // c5t25i2
	assign leaf[36] = !f[326] && f[296] && f[246] && !f[357]; // c5t25i2
	assign leaf[37] = !f[326] && f[296] && f[246] && f[357]; // c5t25i2
	assign leaf[38] = f[326] && !f[304] && !f[322] && !f[332]; // c5t25i2
	assign leaf[39] = f[326] && !f[304] && !f[322] && f[332]; // c5t25i2
	assign leaf[40] = f[326] && !f[304] && f[322] && !f[298]; // c5t25i2
	assign leaf[41] = f[326] && !f[304] && f[322] && f[298]; // c5t25i2
	assign leaf[42] = f[326] && f[304] && !f[381] && !f[215]; // c5t25i2
	assign leaf[43] = f[326] && f[304] && !f[381] && f[215]; // c5t25i2
	assign leaf[44] = f[326] && f[304] && f[381] && !f[322]; // c5t25i2
	assign leaf[45] = f[326] && f[304] && f[381] && f[322]; // c5t25i2
	assign leaf[46] = !f[489] && !f[298] && !f[300] && !f[295]; // c5t35i3
	assign leaf[47] = !f[489] && !f[298] && !f[300] && f[295]; // c5t35i3
	assign leaf[48] = !f[489] && !f[298] && f[300] && !f[328]; // c5t35i3
	assign leaf[49] = !f[489] && !f[298] && f[300] && f[328]; // c5t35i3
	assign leaf[50] = !f[489] && f[298] && !f[275] && !f[219]; // c5t35i3
	assign leaf[51] = !f[489] && f[298] && !f[275] && f[219]; // c5t35i3
	assign leaf[52] = !f[489] && f[298] && f[275] && !f[357]; // c5t35i3
	assign leaf[53] = !f[489] && f[298] && f[275] && f[357]; // c5t35i3
	assign leaf[54] = f[489] && !f[248] && !f[407] && !f[437]; // c5t35i3
	assign leaf[55] = f[489] && !f[248] && !f[407] && f[437]; // c5t35i3
	assign leaf[56] = f[489] && !f[248] && f[407] && !f[276]; // c5t35i3
	assign leaf[57] = f[489] && !f[248] && f[407] && f[276]; // c5t35i3
	assign leaf[58] = f[489] && f[248] && !f[355] && !f[385]; // c5t35i3
	assign leaf[59] = f[489] && f[248] && !f[355] && f[385]; // c5t35i3
	assign leaf[60] = f[489] && f[248] && f[355] && !f[323]; // c5t35i3
	assign leaf[61] = f[489] && f[248] && f[355] && f[323]; // c5t35i3
	assign leaf[62] = !f[375] && !f[320] && !f[191] && !f[248]; // c5t45i4
	assign leaf[63] = !f[375] && !f[320] && !f[191] && f[248]; // c5t45i4
	assign leaf[64] = !f[375] && !f[320] && f[191] && !f[300]; // c5t45i4
	assign leaf[65] = !f[375] && !f[320] && f[191] && f[300]; // c5t45i4
	assign leaf[66] = !f[375] && f[320] && !f[434] && !f[267]; // c5t45i4
	assign leaf[67] = !f[375] && f[320] && !f[434] && f[267]; // c5t45i4
	assign leaf[68] = !f[375] && f[320] && f[434] && !f[380]; // c5t45i4
	assign leaf[69] = !f[375] && f[320] && f[434] && f[380]; // c5t45i4
	assign leaf[70] = f[375] && !f[486] && !f[297] && !f[299]; // c5t45i4
	assign leaf[71] = f[375] && !f[486] && !f[297] && f[299]; // c5t45i4
	assign leaf[72] = f[375] && !f[486] && f[297] && !f[274]; // c5t45i4
	assign leaf[73] = f[375] && !f[486] && f[297] && f[274]; // c5t45i4
	assign leaf[74] = f[375] && f[486] && !f[514] && !f[484]; // c5t45i4
	assign leaf[75] = f[375] && f[486] && !f[514] && f[484]; // c5t45i4
	assign leaf[76] = f[375] && f[486] && f[514] && !f[458]; // c5t45i4
	assign leaf[77] = f[375] && f[486] && f[514] && f[458]; // c5t45i4
	assign leaf[78] = !f[327] && !f[296] && !f[517] && !f[330]; // c5t55i5
	assign leaf[79] = !f[327] && !f[296] && !f[517] && f[330]; // c5t55i5
	assign leaf[80] = !f[327] && !f[296] && f[517] && !f[217]; // c5t55i5
	assign leaf[81] = !f[327] && !f[296] && f[517] && f[217]; // c5t55i5
	assign leaf[82] = !f[327] && f[296] && !f[273] && !f[218]; // c5t55i5
	assign leaf[83] = !f[327] && f[296] && !f[273] && f[218]; // c5t55i5
	assign leaf[84] = !f[327] && f[296] && f[273] && !f[358]; // c5t55i5
	assign leaf[85] = !f[327] && f[296] && f[273] && f[358]; // c5t55i5
	assign leaf[86] = f[327] && !f[323] && !f[305] && !f[382]; // c5t55i5
	assign leaf[87] = f[327] && !f[323] && !f[305] && f[382]; // c5t55i5
	assign leaf[88] = f[327] && !f[323] && f[305] && !f[381]; // c5t55i5
	assign leaf[89] = f[327] && !f[323] && f[305] && f[381]; // c5t55i5
	assign leaf[90] = f[327] && f[323] && !f[409] && !f[522]; // c5t55i5
	assign leaf[91] = f[327] && f[323] && !f[409] && f[522]; // c5t55i5
	assign leaf[92] = f[327] && f[323] && f[409] && !f[248]; // c5t55i5
	assign leaf[93] = f[327] && f[323] && f[409] && f[248]; // c5t55i5
	assign leaf[94] = !f[489] && !f[298] && !f[267] && !f[301]; // c5t65i6
	assign leaf[95] = !f[489] && !f[298] && !f[267] && f[301]; // c5t65i6
	assign leaf[96] = !f[489] && !f[298] && f[267] && !f[243]; // c5t65i6
	assign leaf[97] = !f[489] && !f[298] && f[267] && f[243]; // c5t65i6
	assign leaf[98] = !f[489] && f[298] && !f[275] && !f[304]; // c5t65i6
	assign leaf[99] = !f[489] && f[298] && !f[275] && f[304]; // c5t65i6
	assign leaf[100] = !f[489] && f[298] && f[275] && !f[186]; // c5t65i6
	assign leaf[101] = !f[489] && f[298] && f[275] && f[186]; // c5t65i6
	assign leaf[102] = f[489] && !f[380] && !f[410] && !f[378]; // c5t65i6
	assign leaf[103] = f[489] && !f[380] && !f[410] && f[378]; // c5t65i6
	assign leaf[104] = f[489] && !f[380] && f[410] && !f[352]; // c5t65i6
	assign leaf[105] = f[489] && !f[380] && f[410] && f[352]; // c5t65i6
	assign leaf[106] = f[489] && f[380] && !f[510] && !f[537]; // c5t65i6
	assign leaf[107] = f[489] && f[380] && !f[510] && f[537]; // c5t65i6
	assign leaf[108] = f[489] && f[380] && f[510] && !f[461]; // c5t65i6
	assign leaf[109] = f[489] && f[380] && f[510] && f[461]; // c5t65i6
	assign leaf[110] = !f[490] && !f[297] && !f[300] && !f[186]; // c5t75i7
	assign leaf[111] = !f[490] && !f[297] && !f[300] && f[186]; // c5t75i7
	assign leaf[112] = !f[490] && !f[297] && f[300] && !f[328]; // c5t75i7
	assign leaf[113] = !f[490] && !f[297] && f[300] && f[328]; // c5t75i7
	assign leaf[114] = !f[490] && f[297] && !f[294] && !f[277]; // c5t75i7
	assign leaf[115] = !f[490] && f[297] && !f[294] && f[277]; // c5t75i7
	assign leaf[116] = !f[490] && f[297] && f[294] && !f[241]; // c5t75i7
	assign leaf[117] = !f[490] && f[297] && f[294] && f[241]; // c5t75i7
	assign leaf[118] = f[490] && !f[381] && !f[245] && !f[379]; // c5t75i7
	assign leaf[119] = f[490] && !f[381] && !f[245] && f[379]; // c5t75i7
	assign leaf[120] = f[490] && !f[381] && f[245] && !f[384]; // c5t75i7
	assign leaf[121] = f[490] && !f[381] && f[245] && f[384]; // c5t75i7
	assign leaf[122] = f[490] && f[381] && !f[435] && !f[510]; // c5t75i7
	assign leaf[123] = f[490] && f[381] && !f[435] && f[510]; // c5t75i7
	assign leaf[124] = f[490] && f[381] && f[435] && !f[221]; // c5t75i7
	assign leaf[125] = f[490] && f[381] && f[435] && f[221]; // c5t75i7
	assign leaf[126] = !f[488] && !f[188] && !f[247] && !f[158]; // c5t85i8
	assign leaf[127] = !f[488] && !f[188] && !f[247] && f[158]; // c5t85i8
	assign leaf[128] = !f[488] && !f[188] && f[247] && !f[356]; // c5t85i8
	assign leaf[129] = !f[488] && !f[188] && f[247] && f[356]; // c5t85i8
	assign leaf[130] = !f[488] && f[188] && !f[272] && !f[303]; // c5t85i8
	assign leaf[131] = !f[488] && f[188] && !f[272] && f[303]; // c5t85i8
	assign leaf[132] = !f[488] && f[188] && f[272] && !f[219]; // c5t85i8
	assign leaf[133] = !f[488] && f[188] && f[272] && f[219]; // c5t85i8
	assign leaf[134] = f[488] && !f[380] && !f[410] && !f[374]; // c5t85i8
	assign leaf[135] = f[488] && !f[380] && !f[410] && f[374]; // c5t85i8
	assign leaf[136] = f[488] && !f[380] && f[410] && !f[583]; // c5t85i8
	assign leaf[137] = f[488] && !f[380] && f[410] && f[583]; // c5t85i8
	assign leaf[138] = f[488] && f[380] && !f[461] && !f[245]; // c5t85i8
	assign leaf[139] = f[488] && f[380] && !f[461] && f[245]; // c5t85i8
	assign leaf[140] = f[488] && f[380] && f[461] && !f[353]; // c5t85i8
	assign leaf[141] = f[488] && f[380] && f[461] && f[353]; // c5t85i8
	assign leaf[142] = !f[463] && !f[269] && !f[266] && !f[271]; // c5t95i9
	assign leaf[143] = !f[463] && !f[269] && !f[266] && f[271]; // c5t95i9
	assign leaf[144] = !f[463] && !f[269] && f[266] && !f[215]; // c5t95i9
	assign leaf[145] = !f[463] && !f[269] && f[266] && f[215]; // c5t95i9
	assign leaf[146] = !f[463] && f[269] && !f[245] && !f[305]; // c5t95i9
	assign leaf[147] = !f[463] && f[269] && !f[245] && f[305]; // c5t95i9
	assign leaf[148] = !f[463] && f[269] && f[245] && !f[386]; // c5t95i9
	assign leaf[149] = !f[463] && f[269] && f[245] && f[386]; // c5t95i9
	assign leaf[150] = f[463] && !f[353] && !f[383] && !f[351]; // c5t95i9
	assign leaf[151] = f[463] && !f[353] && !f[383] && f[351]; // c5t95i9
	assign leaf[152] = f[463] && !f[353] && f[383] && !f[525]; // c5t95i9
	assign leaf[153] = f[463] && !f[353] && f[383] && f[525]; // c5t95i9
	assign leaf[154] = f[463] && f[353] && !f[304] && !f[322]; // c5t95i9
	assign leaf[155] = f[463] && f[353] && !f[304] && f[322]; // c5t95i9
	assign leaf[156] = f[463] && f[353] && f[304] && !f[213]; // c5t95i9
	assign leaf[157] = f[463] && f[353] && f[304] && f[213]; // c5t95i9
	assign leaf[158] = !f[487] && !f[598] && !f[546] && !f[296]; // c5t105i10
	assign leaf[159] = !f[487] && !f[598] && !f[546] && f[296]; // c5t105i10
	assign leaf[160] = !f[487] && !f[598] && f[546] && !f[542]; // c5t105i10
	assign leaf[161] = !f[487] && !f[598] && f[546] && f[542]; // c5t105i10
	assign leaf[162] = !f[487] && f[598] && !f[456] && !f[133]; // c5t105i10
	assign leaf[163] = !f[487] && f[598] && !f[456] && f[133]; // c5t105i10
	assign leaf[164] = !f[487] && f[598] && f[456] && !f[484]; // c5t105i10
	assign leaf[165] = !f[487] && f[598] && f[456] && f[484]; // c5t105i10
	assign leaf[166] = f[487] && !f[247] && !f[660] && !f[275]; // c5t105i10
	assign leaf[167] = f[487] && !f[247] && !f[660] && f[275]; // c5t105i10
	assign leaf[168] = f[487] && !f[247] && f[660] && !f[297]; // c5t105i10
	assign leaf[169] = f[487] && !f[247] && f[660] && f[297]; // c5t105i10
	assign leaf[170] = f[487] && f[247] && !f[356] && !f[268]; // c5t105i10
	assign leaf[171] = f[487] && f[247] && !f[356] && f[268]; // c5t105i10
	assign leaf[172] = f[487] && f[247] && f[356] && !f[710]; // c5t105i10
	assign leaf[173] = f[487] && f[247] && f[356] && f[710]; // c5t105i10
	assign leaf[174] = !f[190] && !f[248] && !f[491] && !f[268]; // c5t115i11
	assign leaf[175] = !f[190] && !f[248] && !f[491] && f[268]; // c5t115i11
	assign leaf[176] = !f[190] && !f[248] && f[491] && !f[304]; // c5t115i11
	assign leaf[177] = !f[190] && !f[248] && f[491] && f[304]; // c5t115i11
	assign leaf[178] = !f[190] && f[248] && !f[355] && !f[359]; // c5t115i11
	assign leaf[179] = !f[190] && f[248] && !f[355] && f[359]; // c5t115i11
	assign leaf[180] = !f[190] && f[248] && f[355] && !f[350]; // c5t115i11
	assign leaf[181] = !f[190] && f[248] && f[355] && f[350]; // c5t115i11
	assign leaf[182] = f[190] && !f[301] && !f[303] && !f[299]; // c5t115i11
	assign leaf[183] = f[190] && !f[301] && !f[303] && f[299]; // c5t115i11
	assign leaf[184] = f[190] && !f[301] && f[303] && !f[434]; // c5t115i11
	assign leaf[185] = f[190] && !f[301] && f[303] && f[434]; // c5t115i11
	assign leaf[186] = f[190] && f[301] && !f[269]; // c5t115i11
	assign leaf[187] = f[190] && f[301] && f[269] && !f[329]; // c5t115i11
	assign leaf[188] = f[190] && f[301] && f[269] && f[329]; // c5t115i11
	assign leaf[189] = !f[485] && !f[160] && !f[218] && !f[435]; // c5t125i12
	assign leaf[190] = !f[485] && !f[160] && !f[218] && f[435]; // c5t125i12
	assign leaf[191] = !f[485] && !f[160] && f[218] && !f[331]; // c5t125i12
	assign leaf[192] = !f[485] && !f[160] && f[218] && f[331]; // c5t125i12
	assign leaf[193] = !f[485] && f[160] && !f[271] && !f[246]; // c5t125i12
	assign leaf[194] = !f[485] && f[160] && !f[271] && f[246]; // c5t125i12
	assign leaf[195] = !f[485] && f[160] && f[271] && !f[687]; // c5t125i12
	assign leaf[196] = !f[485] && f[160] && f[271] && f[687]; // c5t125i12
	assign leaf[197] = f[485] && !f[458] && !f[428] && !f[349]; // c5t125i12
	assign leaf[198] = f[485] && !f[458] && !f[428] && f[349]; // c5t125i12
	assign leaf[199] = f[485] && !f[458] && f[428] && !f[512]; // c5t125i12
	assign leaf[200] = f[485] && !f[458] && f[428] && f[512]; // c5t125i12
	assign leaf[201] = f[485] && f[458] && !f[513] && !f[355]; // c5t125i12
	assign leaf[202] = f[485] && f[458] && !f[513] && f[355]; // c5t125i12
	assign leaf[203] = f[485] && f[458] && f[513] && !f[177]; // c5t125i12
	assign leaf[204] = f[485] && f[458] && f[513] && f[177]; // c5t125i12
	assign leaf[205] = !f[346] && !f[459] && !f[568] && !f[189]; // c5t135i13
	assign leaf[206] = !f[346] && !f[459] && !f[568] && f[189]; // c5t135i13
	assign leaf[207] = !f[346] && !f[459] && f[568] && !f[293]; // c5t135i13
	assign leaf[208] = !f[346] && !f[459] && f[568] && f[293]; // c5t135i13
	assign leaf[209] = !f[346] && f[459] && !f[276] && !f[325]; // c5t135i13
	assign leaf[210] = !f[346] && f[459] && !f[276] && f[325]; // c5t135i13
	assign leaf[211] = !f[346] && f[459] && f[276] && !f[380]; // c5t135i13
	assign leaf[212] = !f[346] && f[459] && f[276] && f[380]; // c5t135i13
	assign leaf[213] = f[346] && !f[206] && !f[381] && !f[439]; // c5t135i13
	assign leaf[214] = f[346] && !f[206] && !f[381] && f[439]; // c5t135i13
	assign leaf[215] = f[346] && !f[206] && f[381] && !f[463]; // c5t135i13
	assign leaf[216] = f[346] && !f[206] && f[381] && f[463]; // c5t135i13
	assign leaf[217] = f[346] && f[206] && !f[269] && !f[266]; // c5t135i13
	assign leaf[218] = f[346] && f[206] && !f[269] && f[266]; // c5t135i13
	assign leaf[219] = f[346] && f[206] && f[269] && !f[238]; // c5t135i13
	assign leaf[220] = f[346] && f[206] && f[269] && f[238]; // c5t135i13
	assign leaf[221] = !f[488] && !f[457] && !f[159] && !f[217]; // c5t145i14
	assign leaf[222] = !f[488] && !f[457] && !f[159] && f[217]; // c5t145i14
	assign leaf[223] = !f[488] && !f[457] && f[159] && !f[271]; // c5t145i14
	assign leaf[224] = !f[488] && !f[457] && f[159] && f[271]; // c5t145i14
	assign leaf[225] = !f[488] && f[457] && !f[513] && !f[483]; // c5t145i14
	assign leaf[226] = !f[488] && f[457] && !f[513] && f[483]; // c5t145i14
	assign leaf[227] = !f[488] && f[457] && f[513] && !f[430]; // c5t145i14
	assign leaf[228] = !f[488] && f[457] && f[513] && f[430]; // c5t145i14
	assign leaf[229] = f[488] && !f[380] && !f[686] && !f[276]; // c5t145i14
	assign leaf[230] = f[488] && !f[380] && !f[686] && f[276]; // c5t145i14
	assign leaf[231] = f[488] && !f[380] && f[686] && !f[378]; // c5t145i14
	assign leaf[232] = f[488] && !f[380] && f[686] && f[378]; // c5t145i14
	assign leaf[233] = f[488] && f[380] && !f[434] && !f[540]; // c5t145i14
	assign leaf[234] = f[488] && f[380] && !f[434] && f[540]; // c5t145i14
	assign leaf[235] = f[488] && f[380] && f[434] && !f[551]; // c5t145i14
	assign leaf[236] = f[488] && f[380] && f[434] && f[551]; // c5t145i14
	assign leaf[237] = !f[490] && !f[235] && !f[247] && !f[261]; // c5t155i15
	assign leaf[238] = !f[490] && !f[235] && !f[247] && f[261]; // c5t155i15
	assign leaf[239] = !f[490] && !f[235] && f[247] && !f[387]; // c5t155i15
	assign leaf[240] = !f[490] && !f[235] && f[247] && f[387]; // c5t155i15
	assign leaf[241] = !f[490] && f[235] && !f[299] && !f[330]; // c5t155i15
	assign leaf[242] = !f[490] && f[235] && !f[299] && f[330]; // c5t155i15
	assign leaf[243] = !f[490] && f[235] && f[299] && !f[294]; // c5t155i15
	assign leaf[244] = !f[490] && f[235] && f[299] && f[294]; // c5t155i15
	assign leaf[245] = f[490] && !f[380] && !f[438] && !f[350]; // c5t155i15
	assign leaf[246] = f[490] && !f[380] && !f[438] && f[350]; // c5t155i15
	assign leaf[247] = f[490] && !f[380] && f[438] && !f[686]; // c5t155i15
	assign leaf[248] = f[490] && !f[380] && f[438] && f[686]; // c5t155i15
	assign leaf[249] = f[490] && f[380] && !f[538] && !f[247]; // c5t155i15
	assign leaf[250] = f[490] && f[380] && !f[538] && f[247]; // c5t155i15
	assign leaf[251] = f[490] && f[380] && f[538] && !f[354]; // c5t155i15
	assign leaf[252] = f[490] && f[380] && f[538] && f[354]; // c5t155i15
	assign leaf[253] = !f[435] && !f[493] && !f[289] && !f[379]; // c5t165i16
	assign leaf[254] = !f[435] && !f[493] && !f[289] && f[379]; // c5t165i16
	assign leaf[255] = !f[435] && !f[493] && f[289] && !f[387]; // c5t165i16
	assign leaf[256] = !f[435] && !f[493] && f[289] && f[387]; // c5t165i16
	assign leaf[257] = !f[435] && f[493] && !f[328] && !f[216]; // c5t165i16
	assign leaf[258] = !f[435] && f[493] && !f[328] && f[216]; // c5t165i16
	assign leaf[259] = !f[435] && f[493] && f[328] && !f[133]; // c5t165i16
	assign leaf[260] = !f[435] && f[493] && f[328] && f[133]; // c5t165i16
	assign leaf[261] = f[435] && !f[353] && !f[383] && !f[323]; // c5t165i16
	assign leaf[262] = f[435] && !f[353] && !f[383] && f[323]; // c5t165i16
	assign leaf[263] = f[435] && !f[353] && f[383] && !f[468]; // c5t165i16
	assign leaf[264] = f[435] && !f[353] && f[383] && f[468]; // c5t165i16
	assign leaf[265] = f[435] && f[353] && !f[333] && !f[191]; // c5t165i16
	assign leaf[266] = f[435] && f[353] && !f[333] && f[191]; // c5t165i16
	assign leaf[267] = f[435] && f[353] && f[333]; // c5t165i16
	assign leaf[268] = !f[435] && !f[464] && !f[455] && !f[289]; // c5t175i17
	assign leaf[269] = !f[435] && !f[464] && !f[455] && f[289]; // c5t175i17
	assign leaf[270] = !f[435] && !f[464] && f[455] && !f[522]; // c5t175i17
	assign leaf[271] = !f[435] && !f[464] && f[455] && f[522]; // c5t175i17
	assign leaf[272] = !f[435] && f[464] && !f[383] && !f[468]; // c5t175i17
	assign leaf[273] = !f[435] && f[464] && !f[383] && f[468]; // c5t175i17
	assign leaf[274] = !f[435] && f[464] && f[383] && !f[509]; // c5t175i17
	assign leaf[275] = !f[435] && f[464] && f[383] && f[509]; // c5t175i17
	assign leaf[276] = f[435] && !f[353] && !f[383] && !f[244]; // c5t175i17
	assign leaf[277] = f[435] && !f[353] && !f[383] && f[244]; // c5t175i17
	assign leaf[278] = f[435] && !f[353] && f[383] && !f[497]; // c5t175i17
	assign leaf[279] = f[435] && !f[353] && f[383] && f[497]; // c5t175i17
	assign leaf[280] = f[435] && f[353] && !f[276] && !f[191]; // c5t175i17
	assign leaf[281] = f[435] && f[353] && !f[276] && f[191]; // c5t175i17
	assign leaf[282] = f[435] && f[353] && f[276] && !f[324]; // c5t175i17
	assign leaf[283] = f[435] && f[353] && f[276] && f[324]; // c5t175i17
	assign leaf[284] = !f[277] && !f[461] && !f[130] && !f[187]; // c5t185i18
	assign leaf[285] = !f[277] && !f[461] && !f[130] && f[187]; // c5t185i18
	assign leaf[286] = !f[277] && !f[461] && f[130] && !f[243]; // c5t185i18
	assign leaf[287] = !f[277] && !f[461] && f[130] && f[243]; // c5t185i18
	assign leaf[288] = !f[277] && f[461] && !f[380] && !f[411]; // c5t185i18
	assign leaf[289] = !f[277] && f[461] && !f[380] && f[411]; // c5t185i18
	assign leaf[290] = !f[277] && f[461] && f[380] && !f[325]; // c5t185i18
	assign leaf[291] = !f[277] && f[461] && f[380] && f[325]; // c5t185i18
	assign leaf[292] = f[277] && !f[383] && !f[183] && !f[300]; // c5t185i18
	assign leaf[293] = f[277] && !f[383] && !f[183] && f[300]; // c5t185i18
	assign leaf[294] = f[277] && !f[383] && f[183] && !f[244]; // c5t185i18
	assign leaf[295] = f[277] && !f[383] && f[183] && f[244]; // c5t185i18
	assign leaf[296] = f[277] && f[383]; // c5t185i18
	assign leaf[297] = !f[374] && !f[321] && !f[325] && !f[402]; // c5t195i19
	assign leaf[298] = !f[374] && !f[321] && !f[325] && f[402]; // c5t195i19
	assign leaf[299] = !f[374] && !f[321] && f[325] && !f[380]; // c5t195i19
	assign leaf[300] = !f[374] && !f[321] && f[325] && f[380]; // c5t195i19
	assign leaf[301] = !f[374] && f[321] && !f[568] && !f[187]; // c5t195i19
	assign leaf[302] = !f[374] && f[321] && !f[568] && f[187]; // c5t195i19
	assign leaf[303] = !f[374] && f[321] && f[568] && !f[458]; // c5t195i19
	assign leaf[304] = !f[374] && f[321] && f[568] && f[458]; // c5t195i19
	assign leaf[305] = f[374] && !f[456] && !f[380] && !f[410]; // c5t195i19
	assign leaf[306] = f[374] && !f[456] && !f[380] && f[410]; // c5t195i19
	assign leaf[307] = f[374] && !f[456] && f[380] && !f[463]; // c5t195i19
	assign leaf[308] = f[374] && !f[456] && f[380] && f[463]; // c5t195i19
	assign leaf[309] = f[374] && f[456] && !f[540] && !f[686]; // c5t195i19
	assign leaf[310] = f[374] && f[456] && !f[540] && f[686]; // c5t195i19
	assign leaf[311] = f[374] && f[456] && f[540] && !f[163]; // c5t195i19
	assign leaf[312] = f[374] && f[456] && f[540] && f[163]; // c5t195i19
	assign leaf[313] = !f[374] && !f[292] && !f[356] && !f[325]; // c5t205i20
	assign leaf[314] = !f[374] && !f[292] && !f[356] && f[325]; // c5t205i20
	assign leaf[315] = !f[374] && !f[292] && f[356] && !f[471]; // c5t205i20
	assign leaf[316] = !f[374] && !f[292] && f[356] && f[471]; // c5t205i20
	assign leaf[317] = !f[374] && f[292] && !f[130] && !f[187]; // c5t205i20
	assign leaf[318] = !f[374] && f[292] && !f[130] && f[187]; // c5t205i20
	assign leaf[319] = !f[374] && f[292] && f[130] && !f[459]; // c5t205i20
	assign leaf[320] = !f[374] && f[292] && f[130] && f[459]; // c5t205i20
	assign leaf[321] = f[374] && !f[456] && !f[567] && !f[289]; // c5t205i20
	assign leaf[322] = f[374] && !f[456] && !f[567] && f[289]; // c5t205i20
	assign leaf[323] = f[374] && !f[456] && f[567] && !f[125]; // c5t205i20
	assign leaf[324] = f[374] && !f[456] && f[567] && f[125]; // c5t205i20
	assign leaf[325] = f[374] && f[456] && !f[686] && !f[305]; // c5t205i20
	assign leaf[326] = f[374] && f[456] && !f[686] && f[305]; // c5t205i20
	assign leaf[327] = f[374] && f[456] && f[686] && !f[317]; // c5t205i20
	assign leaf[328] = f[374] && f[456] && f[686] && f[317]; // c5t205i20
	assign leaf[329] = !f[461] && !f[305] && !f[459] && !f[131]; // c5t215i21
	assign leaf[330] = !f[461] && !f[305] && !f[459] && f[131]; // c5t215i21
	assign leaf[331] = !f[461] && !f[305] && f[459] && !f[542]; // c5t215i21
	assign leaf[332] = !f[461] && !f[305] && f[459] && f[542]; // c5t215i21
	assign leaf[333] = !f[461] && f[305] && !f[300]; // c5t215i21
	assign leaf[334] = !f[461] && f[305] && f[300] && !f[239]; // c5t215i21
	assign leaf[335] = !f[461] && f[305] && f[300] && f[239]; // c5t215i21
	assign leaf[336] = f[461] && !f[381] && !f[273] && !f[351]; // c5t215i21
	assign leaf[337] = f[461] && !f[381] && !f[273] && f[351]; // c5t215i21
	assign leaf[338] = f[461] && !f[381] && f[273] && !f[412]; // c5t215i21
	assign leaf[339] = f[461] && !f[381] && f[273] && f[412]; // c5t215i21
	assign leaf[340] = f[461] && f[381] && !f[551] && !f[536]; // c5t215i21
	assign leaf[341] = f[461] && f[381] && !f[551] && f[536]; // c5t215i21
	assign leaf[342] = f[461] && f[381] && f[551] && !f[657]; // c5t215i21
	assign leaf[343] = f[461] && f[381] && f[551] && f[657]; // c5t215i21
	assign leaf[344] = !f[627] && !f[304] && !f[216] && !f[273]; // c5t225i22
	assign leaf[345] = !f[627] && !f[304] && !f[216] && f[273]; // c5t225i22
	assign leaf[346] = !f[627] && !f[304] && f[216] && !f[300]; // c5t225i22
	assign leaf[347] = !f[627] && !f[304] && f[216] && f[300]; // c5t225i22
	assign leaf[348] = !f[627] && f[304] && !f[301] && !f[377]; // c5t225i22
	assign leaf[349] = !f[627] && f[304] && !f[301] && f[377]; // c5t225i22
	assign leaf[350] = !f[627] && f[304] && f[301] && !f[359]; // c5t225i22
	assign leaf[351] = !f[627] && f[304] && f[301] && f[359]; // c5t225i22
	assign leaf[352] = f[627] && !f[513] && !f[517] && !f[236]; // c5t225i22
	assign leaf[353] = f[627] && !f[513] && !f[517] && f[236]; // c5t225i22
	assign leaf[354] = f[627] && !f[513] && f[517] && !f[381]; // c5t225i22
	assign leaf[355] = f[627] && !f[513] && f[517] && f[381]; // c5t225i22
	assign leaf[356] = f[627] && f[513] && !f[458] && !f[602]; // c5t225i22
	assign leaf[357] = f[627] && f[513] && !f[458] && f[602]; // c5t225i22
	assign leaf[358] = f[627] && f[513] && f[458] && !f[177]; // c5t225i22
	assign leaf[359] = f[627] && f[513] && f[458] && f[177]; // c5t225i22
	assign leaf[360] = !f[462] && !f[464] && !f[228] && !f[610]; // c5t235i23
	assign leaf[361] = !f[462] && !f[464] && !f[228] && f[610]; // c5t235i23
	assign leaf[362] = !f[462] && !f[464] && f[228] && !f[691]; // c5t235i23
	assign leaf[363] = !f[462] && !f[464] && f[228] && f[691]; // c5t235i23
	assign leaf[364] = !f[462] && f[464] && !f[353] && !f[411]; // c5t235i23
	assign leaf[365] = !f[462] && f[464] && !f[353] && f[411]; // c5t235i23
	assign leaf[366] = !f[462] && f[464] && f[353] && !f[132]; // c5t235i23
	assign leaf[367] = !f[462] && f[464] && f[353] && f[132]; // c5t235i23
	assign leaf[368] = f[462] && !f[353] && !f[383] && !f[271]; // c5t235i23
	assign leaf[369] = f[462] && !f[353] && !f[383] && f[271]; // c5t235i23
	assign leaf[370] = f[462] && !f[353] && f[383] && !f[660]; // c5t235i23
	assign leaf[371] = f[462] && !f[353] && f[383] && f[660]; // c5t235i23
	assign leaf[372] = f[462] && f[353] && !f[331] && !f[247]; // c5t235i23
	assign leaf[373] = f[462] && f[353] && !f[331] && f[247]; // c5t235i23
	assign leaf[374] = f[462] && f[353] && f[331] && !f[321]; // c5t235i23
	assign leaf[375] = f[462] && f[353] && f[331] && f[321]; // c5t235i23
	assign leaf[376] = !f[380] && !f[325] && !f[411] && !f[242]; // c5t245i24
	assign leaf[377] = !f[380] && !f[325] && !f[411] && f[242]; // c5t245i24
	assign leaf[378] = !f[380] && !f[325] && f[411] && !f[520]; // c5t245i24
	assign leaf[379] = !f[380] && !f[325] && f[411] && f[520]; // c5t245i24
	assign leaf[380] = !f[380] && f[325] && !f[270] && !f[239]; // c5t245i24
	assign leaf[381] = !f[380] && f[325] && !f[270] && f[239]; // c5t245i24
	assign leaf[382] = !f[380] && f[325] && f[270] && !f[294]; // c5t245i24
	assign leaf[383] = !f[380] && f[325] && f[270] && f[294]; // c5t245i24
	assign leaf[384] = f[380] && !f[297] && !f[327] && !f[186]; // c5t245i24
	assign leaf[385] = f[380] && !f[297] && !f[327] && f[186]; // c5t245i24
	assign leaf[386] = f[380] && !f[297] && f[327] && !f[350]; // c5t245i24
	assign leaf[387] = f[380] && !f[297] && f[327] && f[350]; // c5t245i24
	assign leaf[388] = f[380] && f[297] && !f[274] && !f[295]; // c5t245i24
	assign leaf[389] = f[380] && f[297] && !f[274] && f[295]; // c5t245i24
	assign leaf[390] = f[380] && f[297] && f[274] && !f[354]; // c5t245i24
	assign leaf[391] = f[380] && f[297] && f[274] && f[354]; // c5t245i24
	assign leaf[392] = !f[102] && !f[305] && !f[188] && !f[246]; // c5t255i25
	assign leaf[393] = !f[102] && !f[305] && !f[188] && f[246]; // c5t255i25
	assign leaf[394] = !f[102] && !f[305] && f[188] && !f[301]; // c5t255i25
	assign leaf[395] = !f[102] && !f[305] && f[188] && f[301]; // c5t255i25
	assign leaf[396] = !f[102] && f[305] && !f[384] && !f[183]; // c5t255i25
	assign leaf[397] = !f[102] && f[305] && !f[384] && f[183]; // c5t255i25
	assign leaf[398] = !f[102] && f[305] && f[384]; // c5t255i25
	assign leaf[399] = f[102] && !f[207] && !f[324] && !f[571]; // c5t255i25
	assign leaf[400] = f[102] && !f[207] && !f[324] && f[571]; // c5t255i25
	assign leaf[401] = f[102] && !f[207] && f[324] && !f[348]; // c5t255i25
	assign leaf[402] = f[102] && !f[207] && f[324] && f[348]; // c5t255i25
	assign leaf[403] = f[102] && f[207] && !f[372] && !f[264]; // c5t255i25
	assign leaf[404] = f[102] && f[207] && !f[372] && f[264]; // c5t255i25
	assign leaf[405] = f[102] && f[207] && f[372]; // c5t255i25
	assign leaf[406] = !f[485] && !f[541] && !f[379] && !f[409]; // c5t265i26
	assign leaf[407] = !f[485] && !f[541] && !f[379] && f[409]; // c5t265i26
	assign leaf[408] = !f[485] && !f[541] && f[379] && !f[324]; // c5t265i26
	assign leaf[409] = !f[485] && !f[541] && f[379] && f[324]; // c5t265i26
	assign leaf[410] = !f[485] && f[541] && !f[427] && !f[487]; // c5t265i26
	assign leaf[411] = !f[485] && f[541] && !f[427] && f[487]; // c5t265i26
	assign leaf[412] = !f[485] && f[541] && f[427] && !f[354]; // c5t265i26
	assign leaf[413] = !f[485] && f[541] && f[427] && f[354]; // c5t265i26
	assign leaf[414] = f[485] && !f[541] && !f[539] && !f[374]; // c5t265i26
	assign leaf[415] = f[485] && !f[541] && !f[539] && f[374]; // c5t265i26
	assign leaf[416] = f[485] && !f[541] && f[539] && !f[444]; // c5t265i26
	assign leaf[417] = f[485] && !f[541] && f[539] && f[444]; // c5t265i26
	assign leaf[418] = f[485] && f[541] && !f[430] && !f[428]; // c5t265i26
	assign leaf[419] = f[485] && f[541] && !f[430] && f[428]; // c5t265i26
	assign leaf[420] = f[485] && f[541] && f[430] && !f[276]; // c5t265i26
	assign leaf[421] = f[485] && f[541] && f[430] && f[276]; // c5t265i26
	assign leaf[422] = !f[102] && !f[583] && !f[455] && !f[538]; // c5t275i27
	assign leaf[423] = !f[102] && !f[583] && !f[455] && f[538]; // c5t275i27
	assign leaf[424] = !f[102] && !f[583] && f[455] && !f[400]; // c5t275i27
	assign leaf[425] = !f[102] && !f[583] && f[455] && f[400]; // c5t275i27
	assign leaf[426] = !f[102] && f[583] && !f[399] && !f[406]; // c5t275i27
	assign leaf[427] = !f[102] && f[583] && !f[399] && f[406]; // c5t275i27
	assign leaf[428] = !f[102] && f[583] && f[399] && !f[482]; // c5t275i27
	assign leaf[429] = !f[102] && f[583] && f[399] && f[482]; // c5t275i27
	assign leaf[430] = f[102] && !f[352] && !f[159] && !f[211]; // c5t275i27
	assign leaf[431] = f[102] && !f[352] && !f[159] && f[211]; // c5t275i27
	assign leaf[432] = f[102] && !f[352] && f[159] && !f[381]; // c5t275i27
	assign leaf[433] = f[102] && !f[352] && f[159] && f[381]; // c5t275i27
	assign leaf[434] = f[102] && f[352] && !f[243] && !f[320]; // c5t275i27
	assign leaf[435] = f[102] && f[352] && !f[243] && f[320]; // c5t275i27
	assign leaf[436] = f[102] && f[352] && f[243]; // c5t275i27
	assign leaf[437] = !f[380] && !f[454] && !f[465] && !f[378]; // c5t285i28
	assign leaf[438] = !f[380] && !f[454] && !f[465] && f[378]; // c5t285i28
	assign leaf[439] = !f[380] && !f[454] && f[465] && !f[383]; // c5t285i28
	assign leaf[440] = !f[380] && !f[454] && f[465] && f[383]; // c5t285i28
	assign leaf[441] = !f[380] && f[454] && !f[407] && !f[399]; // c5t285i28
	assign leaf[442] = !f[380] && f[454] && !f[407] && f[399]; // c5t285i28
	assign leaf[443] = !f[380] && f[454] && f[407] && !f[440]; // c5t285i28
	assign leaf[444] = !f[380] && f[454] && f[407] && f[440]; // c5t285i28
	assign leaf[445] = f[380] && !f[434] && !f[297] && !f[294]; // c5t285i28
	assign leaf[446] = f[380] && !f[434] && !f[297] && f[294]; // c5t285i28
	assign leaf[447] = f[380] && !f[434] && f[297] && !f[154]; // c5t285i28
	assign leaf[448] = f[380] && !f[434] && f[297] && f[154]; // c5t285i28
	assign leaf[449] = f[380] && f[434] && !f[353] && !f[323]; // c5t285i28
	assign leaf[450] = f[380] && f[434] && !f[353] && f[323]; // c5t285i28
	assign leaf[451] = f[380] && f[434] && f[353] && !f[468]; // c5t285i28
	assign leaf[452] = f[380] && f[434] && f[353] && f[468]; // c5t285i28
	assign leaf[453] = !f[228] && !f[292] && !f[609] && !f[103]; // c5t295i29
	assign leaf[454] = !f[228] && !f[292] && !f[609] && f[103]; // c5t295i29
	assign leaf[455] = !f[228] && !f[292] && f[609] && !f[294]; // c5t295i29
	assign leaf[456] = !f[228] && !f[292] && f[609] && f[294]; // c5t295i29
	assign leaf[457] = !f[228] && f[292] && !f[235] && !f[125]; // c5t295i29
	assign leaf[458] = !f[228] && f[292] && !f[235] && f[125]; // c5t295i29
	assign leaf[459] = !f[228] && f[292] && f[235] && !f[457]; // c5t295i29
	assign leaf[460] = !f[228] && f[292] && f[235] && f[457]; // c5t295i29
	assign leaf[461] = f[228] && !f[172]; // c5t295i29
	assign leaf[462] = f[228] && f[172]; // c5t295i29
	assign leaf[463] = !f[684] && !f[600] && !f[603] && !f[440]; // c5t305i30
	assign leaf[464] = !f[684] && !f[600] && !f[603] && f[440]; // c5t305i30
	assign leaf[465] = !f[684] && !f[600] && f[603] && !f[628]; // c5t305i30
	assign leaf[466] = !f[684] && !f[600] && f[603] && f[628]; // c5t305i30
	assign leaf[467] = !f[684] && f[600] && !f[457] && !f[488]; // c5t305i30
	assign leaf[468] = !f[684] && f[600] && !f[457] && f[488]; // c5t305i30
	assign leaf[469] = !f[684] && f[600] && f[457] && !f[485]; // c5t305i30
	assign leaf[470] = !f[684] && f[600] && f[457] && f[485]; // c5t305i30
	assign leaf[471] = f[684] && !f[289] && !f[296] && !f[263]; // c5t305i30
	assign leaf[472] = f[684] && !f[289] && !f[296] && f[263]; // c5t305i30
	assign leaf[473] = f[684] && !f[289] && f[296] && !f[330]; // c5t305i30
	assign leaf[474] = f[684] && !f[289] && f[296] && f[330]; // c5t305i30
	assign leaf[475] = f[684] && f[289] && !f[578] && !f[373]; // c5t305i30
	assign leaf[476] = f[684] && f[289] && !f[578] && f[373]; // c5t305i30
	assign leaf[477] = f[684] && f[289] && f[578] && !f[401]; // c5t305i30
	assign leaf[478] = f[684] && f[289] && f[578] && f[401]; // c5t305i30
	assign leaf[479] = !f[277] && !f[628] && !f[548] && !f[332]; // c5t315i31
	assign leaf[480] = !f[277] && !f[628] && !f[548] && f[332]; // c5t315i31
	assign leaf[481] = !f[277] && !f[628] && f[548] && !f[683]; // c5t315i31
	assign leaf[482] = !f[277] && !f[628] && f[548] && f[683]; // c5t315i31
	assign leaf[483] = !f[277] && f[628] && !f[483] && !f[235]; // c5t315i31
	assign leaf[484] = !f[277] && f[628] && !f[483] && f[235]; // c5t315i31
	assign leaf[485] = !f[277] && f[628] && f[483] && !f[400]; // c5t315i31
	assign leaf[486] = !f[277] && f[628] && f[483] && f[400]; // c5t315i31
	assign leaf[487] = f[277] && !f[274]; // c5t315i31
	assign leaf[488] = f[277] && f[274] && !f[651]; // c5t315i31
	assign leaf[489] = f[277] && f[274] && f[651]; // c5t315i31
	assign leaf[490] = !f[490] && !f[103] && !f[609] && !f[263]; // c5t325i32
	assign leaf[491] = !f[490] && !f[103] && !f[609] && f[263]; // c5t325i32
	assign leaf[492] = !f[490] && !f[103] && f[609] && !f[287]; // c5t325i32
	assign leaf[493] = !f[490] && !f[103] && f[609] && f[287]; // c5t325i32
	assign leaf[494] = !f[490] && f[103] && !f[405] && !f[577]; // c5t325i32
	assign leaf[495] = !f[490] && f[103] && !f[405] && f[577]; // c5t325i32
	assign leaf[496] = !f[490] && f[103] && f[405] && !f[573]; // c5t325i32
	assign leaf[497] = !f[490] && f[103] && f[405] && f[573]; // c5t325i32
	assign leaf[498] = f[490] && !f[304] && !f[354] && !f[324]; // c5t325i32
	assign leaf[499] = f[490] && !f[304] && !f[354] && f[324]; // c5t325i32
	assign leaf[500] = f[490] && !f[304] && f[354] && !f[323]; // c5t325i32
	assign leaf[501] = f[490] && !f[304] && f[354] && f[323]; // c5t325i32
	assign leaf[502] = f[490] && f[304] && !f[300]; // c5t325i32
	assign leaf[503] = f[490] && f[304] && f[300] && !f[599]; // c5t325i32
	assign leaf[504] = f[490] && f[304] && f[300] && f[599]; // c5t325i32
	assign leaf[505] = !f[434] && !f[464] && !f[713] && !f[120]; // c5t335i33
	assign leaf[506] = !f[434] && !f[464] && !f[713] && f[120]; // c5t335i33
	assign leaf[507] = !f[434] && !f[464] && f[713] && !f[465]; // c5t335i33
	assign leaf[508] = !f[434] && !f[464] && f[713] && f[465]; // c5t335i33
	assign leaf[509] = !f[434] && f[464] && !f[350] && !f[377]; // c5t335i33
	assign leaf[510] = !f[434] && f[464] && !f[350] && f[377]; // c5t335i33
	assign leaf[511] = !f[434] && f[464] && f[350] && !f[265]; // c5t335i33
	assign leaf[512] = !f[434] && f[464] && f[350] && f[265]; // c5t335i33
	assign leaf[513] = f[434] && !f[353] && !f[412] && !f[323]; // c5t335i33
	assign leaf[514] = f[434] && !f[353] && !f[412] && f[323]; // c5t335i33
	assign leaf[515] = f[434] && !f[353] && f[412] && !f[500]; // c5t335i33
	assign leaf[516] = f[434] && !f[353] && f[412] && f[500]; // c5t335i33
	assign leaf[517] = f[434] && f[353] && !f[347] && !f[304]; // c5t335i33
	assign leaf[518] = f[434] && f[353] && !f[347] && f[304]; // c5t335i33
	assign leaf[519] = f[434] && f[353] && f[347] && !f[276]; // c5t335i33
	assign leaf[520] = f[434] && f[353] && f[347] && f[276]; // c5t335i33
	assign leaf[521] = !f[228] && !f[191] && !f[248] && !f[269]; // c5t345i34
	assign leaf[522] = !f[228] && !f[191] && !f[248] && f[269]; // c5t345i34
	assign leaf[523] = !f[228] && !f[191] && f[248] && !f[269]; // c5t345i34
	assign leaf[524] = !f[228] && !f[191] && f[248] && f[269]; // c5t345i34
	assign leaf[525] = !f[228] && f[191] && !f[159] && !f[328]; // c5t345i34
	assign leaf[526] = !f[228] && f[191] && !f[159] && f[328]; // c5t345i34
	assign leaf[527] = !f[228] && f[191] && f[159] && !f[248]; // c5t345i34
	assign leaf[528] = !f[228] && f[191] && f[159] && f[248]; // c5t345i34
	assign leaf[529] = f[228] && !f[172]; // c5t345i34
	assign leaf[530] = f[228] && f[172]; // c5t345i34
	assign leaf[531] = !f[188] && !f[245] && !f[240] && !f[157]; // c5t355i35
	assign leaf[532] = !f[188] && !f[245] && !f[240] && f[157]; // c5t355i35
	assign leaf[533] = !f[188] && !f[245] && f[240] && !f[236]; // c5t355i35
	assign leaf[534] = !f[188] && !f[245] && f[240] && f[236]; // c5t355i35
	assign leaf[535] = !f[188] && f[245] && !f[328] && !f[359]; // c5t355i35
	assign leaf[536] = !f[188] && f[245] && !f[328] && f[359]; // c5t355i35
	assign leaf[537] = !f[188] && f[245] && f[328] && !f[276]; // c5t355i35
	assign leaf[538] = !f[188] && f[245] && f[328] && f[276]; // c5t355i35
	assign leaf[539] = f[188] && !f[213] && !f[216] && !f[246]; // c5t355i35
	assign leaf[540] = f[188] && !f[213] && !f[216] && f[246]; // c5t355i35
	assign leaf[541] = f[188] && !f[213] && f[216] && !f[192]; // c5t355i35
	assign leaf[542] = f[188] && !f[213] && f[216] && f[192]; // c5t355i35
	assign leaf[543] = f[188] && f[213] && !f[300] && !f[303]; // c5t355i35
	assign leaf[544] = f[188] && f[213] && !f[300] && f[303]; // c5t355i35
	assign leaf[545] = f[188] && f[213] && f[300] && !f[688]; // c5t355i35
	assign leaf[546] = f[188] && f[213] && f[300] && f[688]; // c5t355i35
	assign leaf[547] = !f[102] && !f[565] && !f[289] && !f[481]; // c5t365i36
	assign leaf[548] = !f[102] && !f[565] && !f[289] && f[481]; // c5t365i36
	assign leaf[549] = !f[102] && !f[565] && f[289] && !f[178]; // c5t365i36
	assign leaf[550] = !f[102] && !f[565] && f[289] && f[178]; // c5t365i36
	assign leaf[551] = !f[102] && f[565] && !f[302] && !f[267]; // c5t365i36
	assign leaf[552] = !f[102] && f[565] && !f[302] && f[267]; // c5t365i36
	assign leaf[553] = !f[102] && f[565] && f[302] && !f[271]; // c5t365i36
	assign leaf[554] = !f[102] && f[565] && f[302] && f[271]; // c5t365i36
	assign leaf[555] = f[102] && !f[242] && !f[324] && !f[206]; // c5t365i36
	assign leaf[556] = f[102] && !f[242] && !f[324] && f[206]; // c5t365i36
	assign leaf[557] = f[102] && !f[242] && f[324] && !f[291]; // c5t365i36
	assign leaf[558] = f[102] && !f[242] && f[324] && f[291]; // c5t365i36
	assign leaf[559] = f[102] && f[242] && !f[347]; // c5t365i36
	assign leaf[560] = f[102] && f[242] && f[347]; // c5t365i36
	assign leaf[561] = !f[333] && !f[485] && !f[160] && !f[218]; // c5t375i37
	assign leaf[562] = !f[333] && !f[485] && !f[160] && f[218]; // c5t375i37
	assign leaf[563] = !f[333] && !f[485] && f[160] && !f[243]; // c5t375i37
	assign leaf[564] = !f[333] && !f[485] && f[160] && f[243]; // c5t375i37
	assign leaf[565] = !f[333] && f[485] && !f[158] && !f[244]; // c5t375i37
	assign leaf[566] = !f[333] && f[485] && !f[158] && f[244]; // c5t375i37
	assign leaf[567] = !f[333] && f[485] && f[158] && !f[577]; // c5t375i37
	assign leaf[568] = !f[333] && f[485] && f[158] && f[577]; // c5t375i37
	assign leaf[569] = f[333] && !f[330]; // c5t375i37
	assign leaf[570] = f[333] && f[330] && !f[571]; // c5t375i37
	assign leaf[571] = f[333] && f[330] && f[571]; // c5t375i37
	assign leaf[572] = !f[103] && !f[380] && !f[455] && !f[539]; // c5t385i38
	assign leaf[573] = !f[103] && !f[380] && !f[455] && f[539]; // c5t385i38
	assign leaf[574] = !f[103] && !f[380] && f[455] && !f[597]; // c5t385i38
	assign leaf[575] = !f[103] && !f[380] && f[455] && f[597]; // c5t385i38
	assign leaf[576] = !f[103] && f[380] && !f[325] && !f[243]; // c5t385i38
	assign leaf[577] = !f[103] && f[380] && !f[325] && f[243]; // c5t385i38
	assign leaf[578] = !f[103] && f[380] && f[325] && !f[321]; // c5t385i38
	assign leaf[579] = !f[103] && f[380] && f[325] && f[321]; // c5t385i38
	assign leaf[580] = f[103] && !f[243] && !f[324] && !f[319]; // c5t385i38
	assign leaf[581] = f[103] && !f[243] && !f[324] && f[319]; // c5t385i38
	assign leaf[582] = f[103] && !f[243] && f[324] && !f[437]; // c5t385i38
	assign leaf[583] = f[103] && !f[243] && f[324] && f[437]; // c5t385i38
	assign leaf[584] = f[103] && f[243]; // c5t385i38
	assign leaf[585] = !f[304] && !f[188] && !f[490] && !f[239]; // c5t395i39
	assign leaf[586] = !f[304] && !f[188] && !f[490] && f[239]; // c5t395i39
	assign leaf[587] = !f[304] && !f[188] && f[490] && !f[273]; // c5t395i39
	assign leaf[588] = !f[304] && !f[188] && f[490] && f[273]; // c5t395i39
	assign leaf[589] = !f[304] && f[188] && !f[212] && !f[216]; // c5t395i39
	assign leaf[590] = !f[304] && f[188] && !f[212] && f[216]; // c5t395i39
	assign leaf[591] = !f[304] && f[188] && f[212] && !f[300]; // c5t395i39
	assign leaf[592] = !f[304] && f[188] && f[212] && f[300]; // c5t395i39
	assign leaf[593] = f[304] && !f[301] && !f[217]; // c5t395i39
	assign leaf[594] = f[304] && !f[301] && f[217]; // c5t395i39
	assign leaf[595] = f[304] && f[301] && !f[383] && !f[234]; // c5t395i39
	assign leaf[596] = f[304] && f[301] && !f[383] && f[234]; // c5t395i39
	assign leaf[597] = f[304] && f[301] && f[383]; // c5t395i39
	assign leaf[598] = !f[276] && !f[200] && !f[332] && !f[329]; // c5t405i40
	assign leaf[599] = !f[276] && !f[200] && !f[332] && f[329]; // c5t405i40
	assign leaf[600] = !f[276] && !f[200] && f[332] && !f[214]; // c5t405i40
	assign leaf[601] = !f[276] && !f[200] && f[332] && f[214]; // c5t405i40
	assign leaf[602] = !f[276] && f[200] && !f[236]; // c5t405i40
	assign leaf[603] = !f[276] && f[200] && f[236]; // c5t405i40
	assign leaf[604] = f[276] && !f[186] && !f[357] && !f[180]; // c5t405i40
	assign leaf[605] = f[276] && !f[186] && !f[357] && f[180]; // c5t405i40
	assign leaf[606] = f[276] && !f[186] && f[357]; // c5t405i40
	assign leaf[607] = f[276] && f[186] && !f[244]; // c5t405i40
	assign leaf[608] = f[276] && f[186] && f[244]; // c5t405i40
	assign leaf[609] = !f[103] && !f[436] && !f[485] && !f[402]; // c5t415i41
	assign leaf[610] = !f[103] && !f[436] && !f[485] && f[402]; // c5t415i41
	assign leaf[611] = !f[103] && !f[436] && f[485] && !f[541]; // c5t415i41
	assign leaf[612] = !f[103] && !f[436] && f[485] && f[541]; // c5t415i41
	assign leaf[613] = !f[103] && f[436] && !f[354] && !f[215]; // c5t415i41
	assign leaf[614] = !f[103] && f[436] && !f[354] && f[215]; // c5t415i41
	assign leaf[615] = !f[103] && f[436] && f[354] && !f[321]; // c5t415i41
	assign leaf[616] = !f[103] && f[436] && f[354] && f[321]; // c5t415i41
	assign leaf[617] = f[103] && !f[245] && !f[576]; // c5t415i41
	assign leaf[618] = f[103] && !f[245] && f[576] && !f[348]; // c5t415i41
	assign leaf[619] = f[103] && !f[245] && f[576] && f[348]; // c5t415i41
	assign leaf[620] = f[103] && f[245]; // c5t415i41
	assign leaf[621] = !f[612] && !f[565] && !f[289] && !f[481]; // c5t425i42
	assign leaf[622] = !f[612] && !f[565] && !f[289] && f[481]; // c5t425i42
	assign leaf[623] = !f[612] && !f[565] && f[289] && !f[205]; // c5t425i42
	assign leaf[624] = !f[612] && !f[565] && f[289] && f[205]; // c5t425i42
	assign leaf[625] = !f[612] && f[565] && !f[454] && !f[294]; // c5t425i42
	assign leaf[626] = !f[612] && f[565] && !f[454] && f[294]; // c5t425i42
	assign leaf[627] = !f[612] && f[565] && f[454] && !f[246]; // c5t425i42
	assign leaf[628] = !f[612] && f[565] && f[454] && f[246]; // c5t425i42
	assign leaf[629] = f[612]; // c5t425i42
	assign leaf[630] = !f[488] && !f[485] && !f[133] && !f[380]; // c5t435i43
	assign leaf[631] = !f[488] && !f[485] && !f[133] && f[380]; // c5t435i43
	assign leaf[632] = !f[488] && !f[485] && f[133] && !f[218]; // c5t435i43
	assign leaf[633] = !f[488] && !f[485] && f[133] && f[218]; // c5t435i43
	assign leaf[634] = !f[488] && f[485] && !f[430] && !f[372]; // c5t435i43
	assign leaf[635] = !f[488] && f[485] && !f[430] && f[372]; // c5t435i43
	assign leaf[636] = !f[488] && f[485] && f[430] && !f[541]; // c5t435i43
	assign leaf[637] = !f[488] && f[485] && f[430] && f[541]; // c5t435i43
	assign leaf[638] = f[488] && !f[717] && !f[430] && !f[183]; // c5t435i43
	assign leaf[639] = f[488] && !f[717] && !f[430] && f[183]; // c5t435i43
	assign leaf[640] = f[488] && !f[717] && f[430] && !f[322]; // c5t435i43
	assign leaf[641] = f[488] && !f[717] && f[430] && f[322]; // c5t435i43
	assign leaf[642] = f[488] && f[717] && !f[632]; // c5t435i43
	assign leaf[643] = f[488] && f[717] && f[632]; // c5t435i43
	assign leaf[644] = !f[411] && !f[301] && !f[217] && !f[295]; // c5t445i44
	assign leaf[645] = !f[411] && !f[301] && !f[217] && f[295]; // c5t445i44
	assign leaf[646] = !f[411] && !f[301] && f[217] && !f[298]; // c5t445i44
	assign leaf[647] = !f[411] && !f[301] && f[217] && f[298]; // c5t445i44
	assign leaf[648] = !f[411] && f[301] && !f[185] && !f[440]; // c5t445i44
	assign leaf[649] = !f[411] && f[301] && !f[185] && f[440]; // c5t445i44
	assign leaf[650] = !f[411] && f[301] && f[185] && !f[269]; // c5t445i44
	assign leaf[651] = !f[411] && f[301] && f[185] && f[269]; // c5t445i44
	assign leaf[652] = f[411] && !f[496] && !f[353] && !f[124]; // c5t445i44
	assign leaf[653] = f[411] && !f[496] && !f[353] && f[124]; // c5t445i44
	assign leaf[654] = f[411] && !f[496] && f[353] && !f[299]; // c5t445i44
	assign leaf[655] = f[411] && !f[496] && f[353] && f[299]; // c5t445i44
	assign leaf[656] = f[411] && f[496] && !f[185] && !f[127]; // c5t445i44
	assign leaf[657] = f[411] && f[496] && !f[185] && f[127]; // c5t445i44
	assign leaf[658] = f[411] && f[496] && f[185] && !f[271]; // c5t445i44
	assign leaf[659] = f[411] && f[496] && f[185] && f[271]; // c5t445i44
	assign leaf[660] = !f[556] && !f[654] && !f[459] && !f[543]; // c5t455i45
	assign leaf[661] = !f[556] && !f[654] && !f[459] && f[543]; // c5t455i45
	assign leaf[662] = !f[556] && !f[654] && f[459] && !f[401]; // c5t455i45
	assign leaf[663] = !f[556] && !f[654] && f[459] && f[401]; // c5t455i45
	assign leaf[664] = !f[556] && f[654] && !f[264] && !f[153]; // c5t455i45
	assign leaf[665] = !f[556] && f[654] && !f[264] && f[153]; // c5t455i45
	assign leaf[666] = !f[556] && f[654] && f[264] && !f[320]; // c5t455i45
	assign leaf[667] = !f[556] && f[654] && f[264] && f[320]; // c5t455i45
	assign leaf[668] = f[556] && !f[372]; // c5t455i45
	assign leaf[669] = f[556] && f[372] && !f[526]; // c5t455i45
	assign leaf[670] = f[556] && f[372] && f[526] && !f[636]; // c5t455i45
	assign leaf[671] = f[556] && f[372] && f[526] && f[636]; // c5t455i45
	assign leaf[672] = !f[433] && !f[347] && !f[293] && !f[547]; // c5t465i46
	assign leaf[673] = !f[433] && !f[347] && !f[293] && f[547]; // c5t465i46
	assign leaf[674] = !f[433] && !f[347] && f[293] && !f[258]; // c5t465i46
	assign leaf[675] = !f[433] && !f[347] && f[293] && f[258]; // c5t465i46
	assign leaf[676] = !f[433] && f[347] && !f[315] && !f[175]; // c5t465i46
	assign leaf[677] = !f[433] && f[347] && !f[315] && f[175]; // c5t465i46
	assign leaf[678] = !f[433] && f[347] && f[315] && !f[483]; // c5t465i46
	assign leaf[679] = !f[433] && f[347] && f[315] && f[483]; // c5t465i46
	assign leaf[680] = f[433] && !f[352] && !f[382] && !f[385]; // c5t465i46
	assign leaf[681] = f[433] && !f[352] && !f[382] && f[385]; // c5t465i46
	assign leaf[682] = f[433] && !f[352] && f[382] && !f[606]; // c5t465i46
	assign leaf[683] = f[433] && !f[352] && f[382] && f[606]; // c5t465i46
	assign leaf[684] = f[433] && f[352] && !f[331] && !f[468]; // c5t465i46
	assign leaf[685] = f[433] && f[352] && !f[331] && f[468]; // c5t465i46
	assign leaf[686] = f[433] && f[352] && f[331] && !f[275]; // c5t465i46
	assign leaf[687] = f[433] && f[352] && f[331] && f[275]; // c5t465i46
	assign leaf[688] = !f[517] && !f[262] && !f[551] && !f[571]; // c5t475i47
	assign leaf[689] = !f[517] && !f[262] && !f[551] && f[571]; // c5t475i47
	assign leaf[690] = !f[517] && !f[262] && f[551] && !f[236]; // c5t475i47
	assign leaf[691] = !f[517] && !f[262] && f[551] && f[236]; // c5t475i47
	assign leaf[692] = !f[517] && f[262] && !f[178] && !f[351]; // c5t475i47
	assign leaf[693] = !f[517] && f[262] && !f[178] && f[351]; // c5t475i47
	assign leaf[694] = !f[517] && f[262] && f[178] && !f[547]; // c5t475i47
	assign leaf[695] = !f[517] && f[262] && f[178] && f[547]; // c5t475i47
	assign leaf[696] = f[517] && !f[467] && !f[381] && !f[184]; // c5t475i47
	assign leaf[697] = f[517] && !f[467] && !f[381] && f[184]; // c5t475i47
	assign leaf[698] = f[517] && !f[467] && f[381] && !f[513]; // c5t475i47
	assign leaf[699] = f[517] && !f[467] && f[381] && f[513]; // c5t475i47
	assign leaf[700] = f[517] && f[467] && !f[540] && !f[663]; // c5t475i47
	assign leaf[701] = f[517] && f[467] && !f[540] && f[663]; // c5t475i47
	assign leaf[702] = f[517] && f[467] && f[540] && !f[381]; // c5t475i47
	assign leaf[703] = f[517] && f[467] && f[540] && f[381]; // c5t475i47
	assign leaf[704] = !f[264] && !f[241] && !f[239] && !f[243]; // c5t485i48
	assign leaf[705] = !f[264] && !f[241] && !f[239] && f[243]; // c5t485i48
	assign leaf[706] = !f[264] && !f[241] && f[239] && !f[187]; // c5t485i48
	assign leaf[707] = !f[264] && !f[241] && f[239] && f[187]; // c5t485i48
	assign leaf[708] = !f[264] && f[241] && !f[217] && !f[238]; // c5t485i48
	assign leaf[709] = !f[264] && f[241] && !f[217] && f[238]; // c5t485i48
	assign leaf[710] = !f[264] && f[241] && f[217] && !f[239]; // c5t485i48
	assign leaf[711] = !f[264] && f[241] && f[217] && f[239]; // c5t485i48
	assign leaf[712] = f[264] && !f[241] && !f[157] && !f[296]; // c5t485i48
	assign leaf[713] = f[264] && !f[241] && !f[157] && f[296]; // c5t485i48
	assign leaf[714] = f[264] && !f[241] && f[157] && !f[244]; // c5t485i48
	assign leaf[715] = f[264] && !f[241] && f[157] && f[244]; // c5t485i48
	assign leaf[716] = f[264] && f[241] && !f[352] && !f[543]; // c5t485i48
	assign leaf[717] = f[264] && f[241] && !f[352] && f[543]; // c5t485i48
	assign leaf[718] = f[264] && f[241] && f[352] && !f[243]; // c5t485i48
	assign leaf[719] = f[264] && f[241] && f[352] && f[243]; // c5t485i48
	assign leaf[720] = !f[411] && !f[329] && !f[325] && !f[215]; // c5t495i49
	assign leaf[721] = !f[411] && !f[329] && !f[325] && f[215]; // c5t495i49
	assign leaf[722] = !f[411] && !f[329] && f[325] && !f[352]; // c5t495i49
	assign leaf[723] = !f[411] && !f[329] && f[325] && f[352]; // c5t495i49
	assign leaf[724] = !f[411] && f[329] && !f[245] && !f[440]; // c5t495i49
	assign leaf[725] = !f[411] && f[329] && !f[245] && f[440]; // c5t495i49
	assign leaf[726] = !f[411] && f[329] && f[245] && !f[247]; // c5t495i49
	assign leaf[727] = !f[411] && f[329] && f[245] && f[247]; // c5t495i49
	assign leaf[728] = f[411] && !f[329] && !f[179] && !f[237]; // c5t495i49
	assign leaf[729] = f[411] && !f[329] && !f[179] && f[237]; // c5t495i49
	assign leaf[730] = f[411] && !f[329] && f[179] && !f[130]; // c5t495i49
	assign leaf[731] = f[411] && !f[329] && f[179] && f[130]; // c5t495i49
	assign leaf[732] = f[411] && f[329] && !f[150] && !f[130]; // c5t495i49
	assign leaf[733] = f[411] && f[329] && !f[150] && f[130]; // c5t495i49
	assign leaf[734] = f[411] && f[329] && f[150]; // c5t495i49
	assign leaf[735] = !f[102] && !f[556] && !f[433] && !f[468]; // c5t505i50
	assign leaf[736] = !f[102] && !f[556] && !f[433] && f[468]; // c5t505i50
	assign leaf[737] = !f[102] && !f[556] && f[433] && !f[684]; // c5t505i50
	assign leaf[738] = !f[102] && !f[556] && f[433] && f[684]; // c5t505i50
	assign leaf[739] = !f[102] && f[556] && !f[639] && !f[606]; // c5t505i50
	assign leaf[740] = !f[102] && f[556] && !f[639] && f[606]; // c5t505i50
	assign leaf[741] = !f[102] && f[556] && f[639]; // c5t505i50
	assign leaf[742] = f[102] && !f[604] && !f[404]; // c5t505i50
	assign leaf[743] = f[102] && !f[604] && f[404]; // c5t505i50
	assign leaf[744] = f[102] && f[604] && !f[344] && !f[349]; // c5t505i50
	assign leaf[745] = f[102] && f[604] && !f[344] && f[349]; // c5t505i50
	assign leaf[746] = f[102] && f[604] && f[344]; // c5t505i50
	assign leaf[747] = !f[200] && !f[717] && !f[599] && !f[681]; // c5t515i51
	assign leaf[748] = !f[200] && !f[717] && !f[599] && f[681]; // c5t515i51
	assign leaf[749] = !f[200] && !f[717] && f[599] && !f[602]; // c5t515i51
	assign leaf[750] = !f[200] && !f[717] && f[599] && f[602]; // c5t515i51
	assign leaf[751] = !f[200] && f[717] && !f[577] && !f[657]; // c5t515i51
	assign leaf[752] = !f[200] && f[717] && !f[577] && f[657]; // c5t515i51
	assign leaf[753] = !f[200] && f[717] && f[577] && !f[214]; // c5t515i51
	assign leaf[754] = !f[200] && f[717] && f[577] && f[214]; // c5t515i51
	assign leaf[755] = f[200]; // c5t515i51
	assign leaf[756] = !f[264] && !f[241] && !f[243] && !f[239]; // c5t525i52
	assign leaf[757] = !f[264] && !f[241] && !f[243] && f[239]; // c5t525i52
	assign leaf[758] = !f[264] && !f[241] && f[243] && !f[268]; // c5t525i52
	assign leaf[759] = !f[264] && !f[241] && f[243] && f[268]; // c5t525i52
	assign leaf[760] = !f[264] && f[241] && !f[155] && !f[158]; // c5t525i52
	assign leaf[761] = !f[264] && f[241] && !f[155] && f[158]; // c5t525i52
	assign leaf[762] = !f[264] && f[241] && f[155] && !f[238]; // c5t525i52
	assign leaf[763] = !f[264] && f[241] && f[155] && f[238]; // c5t525i52
	assign leaf[764] = f[264] && !f[207] && !f[321] && !f[184]; // c5t525i52
	assign leaf[765] = f[264] && !f[207] && !f[321] && f[184]; // c5t525i52
	assign leaf[766] = f[264] && !f[207] && f[321] && !f[633]; // c5t525i52
	assign leaf[767] = f[264] && !f[207] && f[321] && f[633]; // c5t525i52
	assign leaf[768] = f[264] && f[207] && !f[174] && !f[358]; // c5t525i52
	assign leaf[769] = f[264] && f[207] && !f[174] && f[358]; // c5t525i52
	assign leaf[770] = f[264] && f[207] && f[174] && !f[413]; // c5t525i52
	assign leaf[771] = f[264] && f[207] && f[174] && f[413]; // c5t525i52
	assign leaf[772] = !f[228] && !f[101] && !f[565] && !f[481]; // c5t535i53
	assign leaf[773] = !f[228] && !f[101] && !f[565] && f[481]; // c5t535i53
	assign leaf[774] = !f[228] && !f[101] && f[565] && !f[427]; // c5t535i53
	assign leaf[775] = !f[228] && !f[101] && f[565] && f[427]; // c5t535i53
	assign leaf[776] = !f[228] && f[101] && !f[242] && !f[441]; // c5t535i53
	assign leaf[777] = !f[228] && f[101] && !f[242] && f[441]; // c5t535i53
	assign leaf[778] = !f[228] && f[101] && f[242]; // c5t535i53
	assign leaf[779] = f[228]; // c5t535i53
	assign leaf[780] = !f[382] && !f[440] && !f[324] && !f[270]; // c5t545i54
	assign leaf[781] = !f[382] && !f[440] && !f[324] && f[270]; // c5t545i54
	assign leaf[782] = !f[382] && !f[440] && f[324] && !f[328]; // c5t545i54
	assign leaf[783] = !f[382] && !f[440] && f[324] && f[328]; // c5t545i54
	assign leaf[784] = !f[382] && f[440] && !f[327] && !f[582]; // c5t545i54
	assign leaf[785] = !f[382] && f[440] && !f[327] && f[582]; // c5t545i54
	assign leaf[786] = !f[382] && f[440] && f[327] && !f[272]; // c5t545i54
	assign leaf[787] = !f[382] && f[440] && f[327] && f[272]; // c5t545i54
	assign leaf[788] = f[382] && !f[328] && !f[464] && !f[217]; // c5t545i54
	assign leaf[789] = f[382] && !f[328] && !f[464] && f[217]; // c5t545i54
	assign leaf[790] = f[382] && !f[328] && f[464] && !f[323]; // c5t545i54
	assign leaf[791] = f[382] && !f[328] && f[464] && f[323]; // c5t545i54
	assign leaf[792] = f[382] && f[328] && !f[324] && !f[636]; // c5t545i54
	assign leaf[793] = f[382] && f[328] && !f[324] && f[636]; // c5t545i54
	assign leaf[794] = f[382] && f[328] && f[324] && !f[272]; // c5t545i54
	assign leaf[795] = f[382] && f[328] && f[324] && f[272]; // c5t545i54
	assign leaf[796] = !f[583] && !f[386] && !f[471] && !f[331]; // c5t555i55
	assign leaf[797] = !f[583] && !f[386] && !f[471] && f[331]; // c5t555i55
	assign leaf[798] = !f[583] && !f[386] && f[471] && !f[354]; // c5t555i55
	assign leaf[799] = !f[583] && !f[386] && f[471] && f[354]; // c5t555i55
	assign leaf[800] = !f[583] && f[386] && !f[302] && !f[658]; // c5t555i55
	assign leaf[801] = !f[583] && f[386] && !f[302] && f[658]; // c5t555i55
	assign leaf[802] = !f[583] && f[386] && f[302]; // c5t555i55
	assign leaf[803] = f[583] && !f[230] && !f[176] && !f[398]; // c5t555i55
	assign leaf[804] = f[583] && !f[230] && !f[176] && f[398]; // c5t555i55
	assign leaf[805] = f[583] && !f[230] && f[176] && !f[408]; // c5t555i55
	assign leaf[806] = f[583] && !f[230] && f[176] && f[408]; // c5t555i55
	assign leaf[807] = f[583] && f[230] && !f[287]; // c5t555i55
	assign leaf[808] = f[583] && f[230] && f[287] && !f[238]; // c5t555i55
	assign leaf[809] = f[583] && f[230] && f[287] && f[238]; // c5t555i55
	assign leaf[810] = !f[598] && !f[214] && !f[270] && !f[266]; // c5t565i56
	assign leaf[811] = !f[598] && !f[214] && !f[270] && f[266]; // c5t565i56
	assign leaf[812] = !f[598] && !f[214] && f[270] && !f[294]; // c5t565i56
	assign leaf[813] = !f[598] && !f[214] && f[270] && f[294]; // c5t565i56
	assign leaf[814] = !f[598] && f[214] && !f[297] && !f[327]; // c5t565i56
	assign leaf[815] = !f[598] && f[214] && !f[297] && f[327]; // c5t565i56
	assign leaf[816] = !f[598] && f[214] && f[297] && !f[709]; // c5t565i56
	assign leaf[817] = !f[598] && f[214] && f[297] && f[709]; // c5t565i56
	assign leaf[818] = f[598] && !f[486] && !f[428] && !f[398]; // c5t565i56
	assign leaf[819] = f[598] && !f[486] && !f[428] && f[398]; // c5t565i56
	assign leaf[820] = f[598] && !f[486] && f[428] && !f[483]; // c5t565i56
	assign leaf[821] = f[598] && !f[486] && f[428] && f[483]; // c5t565i56
	assign leaf[822] = f[598] && f[486] && !f[541] && !f[429]; // c5t565i56
	assign leaf[823] = f[598] && f[486] && !f[541] && f[429]; // c5t565i56
	assign leaf[824] = f[598] && f[486] && f[541] && !f[370]; // c5t565i56
	assign leaf[825] = f[598] && f[486] && f[541] && f[370]; // c5t565i56
	assign leaf[826] = !f[129] && !f[215] && !f[273] && !f[239]; // c5t575i57
	assign leaf[827] = !f[129] && !f[215] && !f[273] && f[239]; // c5t575i57
	assign leaf[828] = !f[129] && !f[215] && f[273] && !f[270]; // c5t575i57
	assign leaf[829] = !f[129] && !f[215] && f[273] && f[270]; // c5t575i57
	assign leaf[830] = !f[129] && f[215] && !f[297] && !f[328]; // c5t575i57
	assign leaf[831] = !f[129] && f[215] && !f[297] && f[328]; // c5t575i57
	assign leaf[832] = !f[129] && f[215] && f[297] && !f[293]; // c5t575i57
	assign leaf[833] = !f[129] && f[215] && f[297] && f[293]; // c5t575i57
	assign leaf[834] = f[129] && !f[242] && !f[218] && !f[601]; // c5t575i57
	assign leaf[835] = f[129] && !f[242] && !f[218] && f[601]; // c5t575i57
	assign leaf[836] = f[129] && !f[242] && f[218]; // c5t575i57
	assign leaf[837] = f[129] && f[242] && !f[239]; // c5t575i57
	assign leaf[838] = f[129] && f[242] && f[239] && !f[125]; // c5t575i57
	assign leaf[839] = f[129] && f[242] && f[239] && f[125]; // c5t575i57
	assign leaf[840] = !f[380] && !f[292] && !f[413] && !f[345]; // c5t585i58
	assign leaf[841] = !f[380] && !f[292] && !f[413] && f[345]; // c5t585i58
	assign leaf[842] = !f[380] && !f[292] && f[413] && !f[661]; // c5t585i58
	assign leaf[843] = !f[380] && !f[292] && f[413] && f[661]; // c5t585i58
	assign leaf[844] = !f[380] && f[292] && !f[347] && !f[315]; // c5t585i58
	assign leaf[845] = !f[380] && f[292] && !f[347] && f[315]; // c5t585i58
	assign leaf[846] = !f[380] && f[292] && f[347] && !f[298]; // c5t585i58
	assign leaf[847] = !f[380] && f[292] && f[347] && f[298]; // c5t585i58
	assign leaf[848] = f[380] && !f[131] && !f[349] && !f[659]; // c5t585i58
	assign leaf[849] = f[380] && !f[131] && !f[349] && f[659]; // c5t585i58
	assign leaf[850] = f[380] && !f[131] && f[349] && !f[245]; // c5t585i58
	assign leaf[851] = f[380] && !f[131] && f[349] && f[245]; // c5t585i58
	assign leaf[852] = f[380] && f[131] && !f[630] && !f[550]; // c5t585i58
	assign leaf[853] = f[380] && f[131] && !f[630] && f[550]; // c5t585i58
	assign leaf[854] = f[380] && f[131] && f[630] && !f[651]; // c5t585i58
	assign leaf[855] = f[380] && f[131] && f[630] && f[651]; // c5t585i58
	assign leaf[856] = !f[442] && !f[538] && !f[160] && !f[546]; // c5t595i59
	assign leaf[857] = !f[442] && !f[538] && !f[160] && f[546]; // c5t595i59
	assign leaf[858] = !f[442] && !f[538] && f[160] && !f[513]; // c5t595i59
	assign leaf[859] = !f[442] && !f[538] && f[160] && f[513]; // c5t595i59
	assign leaf[860] = !f[442] && f[538] && !f[400] && !f[316]; // c5t595i59
	assign leaf[861] = !f[442] && f[538] && !f[400] && f[316]; // c5t595i59
	assign leaf[862] = !f[442] && f[538] && f[400] && !f[454]; // c5t595i59
	assign leaf[863] = !f[442] && f[538] && f[400] && f[454]; // c5t595i59
	assign leaf[864] = f[442] && !f[176] && !f[245] && !f[262]; // c5t595i59
	assign leaf[865] = f[442] && !f[176] && !f[245] && f[262]; // c5t595i59
	assign leaf[866] = f[442] && !f[176] && f[245] && !f[567]; // c5t595i59
	assign leaf[867] = f[442] && !f[176] && f[245] && f[567]; // c5t595i59
	assign leaf[868] = f[442] && f[176] && !f[179]; // c5t595i59
	assign leaf[869] = f[442] && f[176] && f[179] && !f[287]; // c5t595i59
	assign leaf[870] = f[442] && f[176] && f[179] && f[287]; // c5t595i59
	assign leaf[871] = !f[713] && !f[630] && !f[403] && !f[511]; // c5t605i60
	assign leaf[872] = !f[713] && !f[630] && !f[403] && f[511]; // c5t605i60
	assign leaf[873] = !f[713] && !f[630] && f[403] && !f[406]; // c5t605i60
	assign leaf[874] = !f[713] && !f[630] && f[403] && f[406]; // c5t605i60
	assign leaf[875] = !f[713] && f[630] && !f[347] && !f[270]; // c5t605i60
	assign leaf[876] = !f[713] && f[630] && !f[347] && f[270]; // c5t605i60
	assign leaf[877] = !f[713] && f[630] && f[347] && !f[263]; // c5t605i60
	assign leaf[878] = !f[713] && f[630] && f[347] && f[263]; // c5t605i60
	assign leaf[879] = f[713] && !f[574] && !f[240] && !f[460]; // c5t605i60
	assign leaf[880] = f[713] && !f[574] && !f[240] && f[460]; // c5t605i60
	assign leaf[881] = f[713] && !f[574] && f[240] && !f[434]; // c5t605i60
	assign leaf[882] = f[713] && !f[574] && f[240] && f[434]; // c5t605i60
	assign leaf[883] = f[713] && f[574] && !f[710] && !f[683]; // c5t605i60
	assign leaf[884] = f[713] && f[574] && !f[710] && f[683]; // c5t605i60
	assign leaf[885] = f[713] && f[574] && f[710]; // c5t605i60
	assign leaf[886] = !f[459] && !f[411] && !f[551] && !f[151]; // c5t615i61
	assign leaf[887] = !f[459] && !f[411] && !f[551] && f[151]; // c5t615i61
	assign leaf[888] = !f[459] && !f[411] && f[551] && !f[294]; // c5t615i61
	assign leaf[889] = !f[459] && !f[411] && f[551] && f[294]; // c5t615i61
	assign leaf[890] = !f[459] && f[411] && !f[329] && !f[179]; // c5t615i61
	assign leaf[891] = !f[459] && f[411] && !f[329] && f[179]; // c5t615i61
	assign leaf[892] = !f[459] && f[411] && f[329]; // c5t615i61
	assign leaf[893] = f[459] && !f[430] && !f[712] && !f[375]; // c5t615i61
	assign leaf[894] = f[459] && !f[430] && !f[712] && f[375]; // c5t615i61
	assign leaf[895] = f[459] && !f[430] && f[712]; // c5t615i61
	assign leaf[896] = f[459] && f[430] && !f[542] && !f[627]; // c5t615i61
	assign leaf[897] = f[459] && f[430] && !f[542] && f[627]; // c5t615i61
	assign leaf[898] = f[459] && f[430] && f[542] && !f[576]; // c5t615i61
	assign leaf[899] = f[459] && f[430] && f[542] && f[576]; // c5t615i61
	assign leaf[900] = !f[402] && !f[630] && !f[270] && !f[126]; // c5t625i62
	assign leaf[901] = !f[402] && !f[630] && !f[270] && f[126]; // c5t625i62
	assign leaf[902] = !f[402] && !f[630] && f[270] && !f[214]; // c5t625i62
	assign leaf[903] = !f[402] && !f[630] && f[270] && f[214]; // c5t625i62
	assign leaf[904] = !f[402] && f[630] && !f[269] && !f[157]; // c5t625i62
	assign leaf[905] = !f[402] && f[630] && !f[269] && f[157]; // c5t625i62
	assign leaf[906] = !f[402] && f[630] && f[269] && !f[265]; // c5t625i62
	assign leaf[907] = !f[402] && f[630] && f[269] && f[265]; // c5t625i62
	assign leaf[908] = f[402] && !f[546] && !f[344] && !f[294]; // c5t625i62
	assign leaf[909] = f[402] && !f[546] && !f[344] && f[294]; // c5t625i62
	assign leaf[910] = f[402] && !f[546] && f[344] && !f[427]; // c5t625i62
	assign leaf[911] = f[402] && !f[546] && f[344] && f[427]; // c5t625i62
	assign leaf[912] = f[402] && f[546] && !f[185] && !f[234]; // c5t625i62
	assign leaf[913] = f[402] && f[546] && !f[185] && f[234]; // c5t625i62
	assign leaf[914] = f[402] && f[546] && f[185] && !f[378]; // c5t625i62
	assign leaf[915] = f[402] && f[546] && f[185] && f[378]; // c5t625i62
	assign leaf[916] = !f[631] && !f[715] && !f[514] && !f[440]; // c5t635i63
	assign leaf[917] = !f[631] && !f[715] && !f[514] && f[440]; // c5t635i63
	assign leaf[918] = !f[631] && !f[715] && f[514] && !f[655]; // c5t635i63
	assign leaf[919] = !f[631] && !f[715] && f[514] && f[655]; // c5t635i63
	assign leaf[920] = !f[631] && f[715] && !f[463] && !f[294]; // c5t635i63
	assign leaf[921] = !f[631] && f[715] && !f[463] && f[294]; // c5t635i63
	assign leaf[922] = !f[631] && f[715] && f[463]; // c5t635i63
	assign leaf[923] = f[631] && !f[457] && !f[159] && !f[553]; // c5t635i63
	assign leaf[924] = f[631] && !f[457] && !f[159] && f[553]; // c5t635i63
	assign leaf[925] = f[631] && !f[457] && f[159] && !f[211]; // c5t635i63
	assign leaf[926] = f[631] && !f[457] && f[159] && f[211]; // c5t635i63
	assign leaf[927] = f[631] && f[457] && !f[712] && !f[398]; // c5t635i63
	assign leaf[928] = f[631] && f[457] && !f[712] && f[398]; // c5t635i63
	assign leaf[929] = f[631] && f[457] && f[712] && !f[295]; // c5t635i63
	assign leaf[930] = f[631] && f[457] && f[712] && f[295]; // c5t635i63
	assign leaf[931] = !f[612] && !f[598] && !f[684] && !f[512]; // c5t645i64
	assign leaf[932] = !f[612] && !f[598] && !f[684] && f[512]; // c5t645i64
	assign leaf[933] = !f[612] && !f[598] && f[684] && !f[576]; // c5t645i64
	assign leaf[934] = !f[612] && !f[598] && f[684] && f[576]; // c5t645i64
	assign leaf[935] = !f[612] && f[598] && !f[486] && !f[428]; // c5t645i64
	assign leaf[936] = !f[612] && f[598] && !f[486] && f[428]; // c5t645i64
	assign leaf[937] = !f[612] && f[598] && f[486] && !f[371]; // c5t645i64
	assign leaf[938] = !f[612] && f[598] && f[486] && f[371]; // c5t645i64
	assign leaf[939] = f[612]; // c5t645i64
	assign leaf[940] = !f[381] && !f[326] && !f[441] && !f[324]; // c5t655i65
	assign leaf[941] = !f[381] && !f[326] && !f[441] && f[324]; // c5t655i65
	assign leaf[942] = !f[381] && !f[326] && f[441] && !f[661]; // c5t655i65
	assign leaf[943] = !f[381] && !f[326] && f[441] && f[661]; // c5t655i65
	assign leaf[944] = !f[381] && f[326] && !f[243] && !f[485]; // c5t655i65
	assign leaf[945] = !f[381] && f[326] && !f[243] && f[485]; // c5t655i65
	assign leaf[946] = !f[381] && f[326] && f[243] && !f[156]; // c5t655i65
	assign leaf[947] = !f[381] && f[326] && f[243] && f[156]; // c5t655i65
	assign leaf[948] = f[381] && !f[327] && !f[132] && !f[244]; // c5t655i65
	assign leaf[949] = f[381] && !f[327] && !f[132] && f[244]; // c5t655i65
	assign leaf[950] = f[381] && !f[327] && f[132] && !f[243]; // c5t655i65
	assign leaf[951] = f[381] && !f[327] && f[132] && f[243]; // c5t655i65
	assign leaf[952] = f[381] && f[327] && !f[294] && !f[409]; // c5t655i65
	assign leaf[953] = f[381] && f[327] && !f[294] && f[409]; // c5t655i65
	assign leaf[954] = f[381] && f[327] && f[294] && !f[653]; // c5t655i65
	assign leaf[955] = f[381] && f[327] && f[294] && f[653]; // c5t655i65
	assign leaf[956] = !f[99] && !f[188] && !f[244] && !f[239]; // c5t665i66
	assign leaf[957] = !f[99] && !f[188] && !f[244] && f[239]; // c5t665i66
	assign leaf[958] = !f[99] && !f[188] && f[244] && !f[267]; // c5t665i66
	assign leaf[959] = !f[99] && !f[188] && f[244] && f[267]; // c5t665i66
	assign leaf[960] = !f[99] && f[188] && !f[273] && !f[271]; // c5t665i66
	assign leaf[961] = !f[99] && f[188] && !f[273] && f[271]; // c5t665i66
	assign leaf[962] = !f[99] && f[188] && f[273] && !f[269]; // c5t665i66
	assign leaf[963] = !f[99] && f[188] && f[273] && f[269]; // c5t665i66
	assign leaf[964] = f[99] && !f[240] && !f[431] && !f[344]; // c5t665i66
	assign leaf[965] = f[99] && !f[240] && !f[431] && f[344]; // c5t665i66
	assign leaf[966] = f[99] && !f[240] && f[431] && !f[317]; // c5t665i66
	assign leaf[967] = f[99] && !f[240] && f[431] && f[317]; // c5t665i66
	assign leaf[968] = f[99] && f[240] && !f[185]; // c5t665i66
	assign leaf[969] = f[99] && f[240] && f[185]; // c5t665i66
	assign leaf[970] = !f[200] && !f[436] && !f[485] && !f[292]; // c5t675i67
	assign leaf[971] = !f[200] && !f[436] && !f[485] && f[292]; // c5t675i67
	assign leaf[972] = !f[200] && !f[436] && f[485] && !f[352]; // c5t675i67
	assign leaf[973] = !f[200] && !f[436] && f[485] && f[352]; // c5t675i67
	assign leaf[974] = !f[200] && f[436] && !f[354] && !f[384]; // c5t675i67
	assign leaf[975] = !f[200] && f[436] && !f[354] && f[384]; // c5t675i67
	assign leaf[976] = !f[200] && f[436] && f[354] && !f[324]; // c5t675i67
	assign leaf[977] = !f[200] && f[436] && f[354] && f[324]; // c5t675i67
	assign leaf[978] = f[200]; // c5t675i67
	assign leaf[979] = !f[120] && !f[686] && !f[598] && !f[509]; // c5t685i68
	assign leaf[980] = !f[120] && !f[686] && !f[598] && f[509]; // c5t685i68
	assign leaf[981] = !f[120] && !f[686] && f[598] && !f[214]; // c5t685i68
	assign leaf[982] = !f[120] && !f[686] && f[598] && f[214]; // c5t685i68
	assign leaf[983] = !f[120] && f[686] && !f[546] && !f[345]; // c5t685i68
	assign leaf[984] = !f[120] && f[686] && !f[546] && f[345]; // c5t685i68
	assign leaf[985] = !f[120] && f[686] && f[546] && !f[682]; // c5t685i68
	assign leaf[986] = !f[120] && f[686] && f[546] && f[682]; // c5t685i68
	assign leaf[987] = f[120] && !f[204] && !f[553]; // c5t685i68
	assign leaf[988] = f[120] && !f[204] && f[553]; // c5t685i68
	assign leaf[989] = f[120] && f[204]; // c5t685i68
	assign leaf[990] = !f[465] && !f[409] && !f[379] && !f[496]; // c5t695i69
	assign leaf[991] = !f[465] && !f[409] && !f[379] && f[496]; // c5t695i69
	assign leaf[992] = !f[465] && !f[409] && f[379] && !f[433]; // c5t695i69
	assign leaf[993] = !f[465] && !f[409] && f[379] && f[433]; // c5t695i69
	assign leaf[994] = !f[465] && f[409] && !f[294] && !f[579]; // c5t695i69
	assign leaf[995] = !f[465] && f[409] && !f[294] && f[579]; // c5t695i69
	assign leaf[996] = !f[465] && f[409] && f[294] && !f[298]; // c5t695i69
	assign leaf[997] = !f[465] && f[409] && f[294] && f[298]; // c5t695i69
	assign leaf[998] = f[465] && !f[355] && !f[296] && !f[376]; // c5t695i69
	assign leaf[999] = f[465] && !f[355] && !f[296] && f[376]; // c5t695i69
	assign leaf[1000] = f[465] && !f[355] && f[296] && !f[301]; // c5t695i69
	assign leaf[1001] = f[465] && !f[355] && f[296] && f[301]; // c5t695i69
	assign leaf[1002] = f[465] && f[355] && !f[509] && !f[624]; // c5t695i69
	assign leaf[1003] = f[465] && f[355] && !f[509] && f[624]; // c5t695i69
	assign leaf[1004] = f[465] && f[355] && f[509] && !f[190]; // c5t695i69
	assign leaf[1005] = f[465] && f[355] && f[509] && f[190]; // c5t695i69
	assign leaf[1006] = !f[120] && !f[630] && !f[714] && !f[270]; // c5t705i70
	assign leaf[1007] = !f[120] && !f[630] && !f[714] && f[270]; // c5t705i70
	assign leaf[1008] = !f[120] && !f[630] && f[714] && !f[296]; // c5t705i70
	assign leaf[1009] = !f[120] && !f[630] && f[714] && f[296]; // c5t705i70
	assign leaf[1010] = !f[120] && f[630] && !f[483] && !f[628]; // c5t705i70
	assign leaf[1011] = !f[120] && f[630] && !f[483] && f[628]; // c5t705i70
	assign leaf[1012] = !f[120] && f[630] && f[483] && !f[345]; // c5t705i70
	assign leaf[1013] = !f[120] && f[630] && f[483] && f[345]; // c5t705i70
	assign leaf[1014] = f[120] && !f[231] && !f[553]; // c5t705i70
	assign leaf[1015] = f[120] && !f[231] && f[553]; // c5t705i70
	assign leaf[1016] = f[120] && f[231]; // c5t705i70
	assign leaf[1017] = !f[382] && !f[440] && !f[301] && !f[324]; // c5t715i71
	assign leaf[1018] = !f[382] && !f[440] && !f[301] && f[324]; // c5t715i71
	assign leaf[1019] = !f[382] && !f[440] && f[301] && !f[186]; // c5t715i71
	assign leaf[1020] = !f[382] && !f[440] && f[301] && f[186]; // c5t715i71
	assign leaf[1021] = !f[382] && f[440] && !f[484] && !f[302]; // c5t715i71
	assign leaf[1022] = !f[382] && f[440] && !f[484] && f[302]; // c5t715i71
	assign leaf[1023] = !f[382] && f[440] && f[484] && !f[383]; // c5t715i71
	assign leaf[1024] = !f[382] && f[440] && f[484] && f[383]; // c5t715i71
	assign leaf[1025] = f[382] && !f[524] && !f[349] && !f[483]; // c5t715i71
	assign leaf[1026] = f[382] && !f[524] && !f[349] && f[483]; // c5t715i71
	assign leaf[1027] = f[382] && !f[524] && f[349] && !f[292]; // c5t715i71
	assign leaf[1028] = f[382] && !f[524] && f[349] && f[292]; // c5t715i71
	assign leaf[1029] = f[382] && f[524] && !f[490] && !f[233]; // c5t715i71
	assign leaf[1030] = f[382] && f[524] && !f[490] && f[233]; // c5t715i71
	assign leaf[1031] = f[382] && f[524] && f[490] && !f[240]; // c5t715i71
	assign leaf[1032] = f[382] && f[524] && f[490] && f[240]; // c5t715i71
	assign leaf[1033] = !f[102] && !f[584] && !f[483] && !f[625]; // c5t725i72
	assign leaf[1034] = !f[102] && !f[584] && !f[483] && f[625]; // c5t725i72
	assign leaf[1035] = !f[102] && !f[584] && f[483] && !f[428]; // c5t725i72
	assign leaf[1036] = !f[102] && !f[584] && f[483] && f[428]; // c5t725i72
	assign leaf[1037] = !f[102] && f[584] && !f[290]; // c5t725i72
	assign leaf[1038] = !f[102] && f[584] && f[290]; // c5t725i72
	assign leaf[1039] = f[102] && !f[603]; // c5t725i72
	assign leaf[1040] = f[102] && f[603] && !f[401] && !f[431]; // c5t725i72
	assign leaf[1041] = f[102] && f[603] && !f[401] && f[431]; // c5t725i72
	assign leaf[1042] = f[102] && f[603] && f[401] && !f[237]; // c5t725i72
	assign leaf[1043] = f[102] && f[603] && f[401] && f[237]; // c5t725i72
	assign leaf[1044] = !f[145] && !f[285] && !f[380] && !f[353]; // c5t735i73
	assign leaf[1045] = !f[145] && !f[285] && !f[380] && f[353]; // c5t735i73
	assign leaf[1046] = !f[145] && !f[285] && f[380] && !f[377]; // c5t735i73
	assign leaf[1047] = !f[145] && !f[285] && f[380] && f[377]; // c5t735i73
	assign leaf[1048] = !f[145] && f[285] && !f[371] && !f[185]; // c5t735i73
	assign leaf[1049] = !f[145] && f[285] && !f[371] && f[185]; // c5t735i73
	assign leaf[1050] = !f[145] && f[285] && f[371] && !f[527]; // c5t735i73
	assign leaf[1051] = !f[145] && f[285] && f[371] && f[527]; // c5t735i73
	assign leaf[1052] = f[145]; // c5t735i73
	assign leaf[1053] = !f[322] && !f[349] && !f[520] && !f[263]; // c5t745i74
	assign leaf[1054] = !f[322] && !f[349] && !f[520] && f[263]; // c5t745i74
	assign leaf[1055] = !f[322] && !f[349] && f[520] && !f[490]; // c5t745i74
	assign leaf[1056] = !f[322] && !f[349] && f[520] && f[490]; // c5t745i74
	assign leaf[1057] = !f[322] && f[349] && !f[174] && !f[267]; // c5t745i74
	assign leaf[1058] = !f[322] && f[349] && !f[174] && f[267]; // c5t745i74
	assign leaf[1059] = !f[322] && f[349] && f[174] && !f[235]; // c5t745i74
	assign leaf[1060] = !f[322] && f[349] && f[174] && f[235]; // c5t745i74
	assign leaf[1061] = f[322] && !f[218] && !f[268] && !f[156]; // c5t745i74
	assign leaf[1062] = f[322] && !f[218] && !f[268] && f[156]; // c5t745i74
	assign leaf[1063] = f[322] && !f[218] && f[268] && !f[295]; // c5t745i74
	assign leaf[1064] = f[322] && !f[218] && f[268] && f[295]; // c5t745i74
	assign leaf[1065] = f[322] && f[218] && !f[160] && !f[273]; // c5t745i74
	assign leaf[1066] = f[322] && f[218] && !f[160] && f[273]; // c5t745i74
	assign leaf[1067] = f[322] && f[218] && f[160] && !f[237]; // c5t745i74
	assign leaf[1068] = f[322] && f[218] && f[160] && f[237]; // c5t745i74
	assign leaf[1069] = !f[402] && !f[484] && !f[631] && !f[493]; // c5t755i75
	assign leaf[1070] = !f[402] && !f[484] && !f[631] && f[493]; // c5t755i75
	assign leaf[1071] = !f[402] && !f[484] && f[631] && !f[601]; // c5t755i75
	assign leaf[1072] = !f[402] && !f[484] && f[631] && f[601]; // c5t755i75
	assign leaf[1073] = !f[402] && f[484] && !f[371] && !f[459]; // c5t755i75
	assign leaf[1074] = !f[402] && f[484] && !f[371] && f[459]; // c5t755i75
	assign leaf[1075] = !f[402] && f[484] && f[371] && !f[430]; // c5t755i75
	assign leaf[1076] = !f[402] && f[484] && f[371] && f[430]; // c5t755i75
	assign leaf[1077] = f[402] && !f[484] && !f[518] && !f[318]; // c5t755i75
	assign leaf[1078] = f[402] && !f[484] && !f[518] && f[318]; // c5t755i75
	assign leaf[1079] = f[402] && !f[484] && f[518] && !f[184]; // c5t755i75
	assign leaf[1080] = f[402] && !f[484] && f[518] && f[184]; // c5t755i75
	assign leaf[1081] = f[402] && f[484] && !f[625] && !f[317]; // c5t755i75
	assign leaf[1082] = f[402] && f[484] && !f[625] && f[317]; // c5t755i75
	assign leaf[1083] = f[402] && f[484] && f[625] && !f[489]; // c5t755i75
	assign leaf[1084] = f[402] && f[484] && f[625] && f[489]; // c5t755i75
	assign leaf[1085] = !f[707] && !f[402] && !f[243] && !f[187]; // c5t765i76
	assign leaf[1086] = !f[707] && !f[402] && !f[243] && f[187]; // c5t765i76
	assign leaf[1087] = !f[707] && !f[402] && f[243] && !f[240]; // c5t765i76
	assign leaf[1088] = !f[707] && !f[402] && f[243] && f[240]; // c5t765i76
	assign leaf[1089] = !f[707] && f[402] && !f[156] && !f[177]; // c5t765i76
	assign leaf[1090] = !f[707] && f[402] && !f[156] && f[177]; // c5t765i76
	assign leaf[1091] = !f[707] && f[402] && f[156] && !f[270]; // c5t765i76
	assign leaf[1092] = !f[707] && f[402] && f[156] && f[270]; // c5t765i76
	assign leaf[1093] = f[707] && !f[627]; // c5t765i76
	assign leaf[1094] = f[707] && f[627]; // c5t765i76
	assign leaf[1095] = !f[190] && !f[130] && !f[406] && !f[464]; // c5t775i77
	assign leaf[1096] = !f[190] && !f[130] && !f[406] && f[464]; // c5t775i77
	assign leaf[1097] = !f[190] && !f[130] && f[406] && !f[325]; // c5t775i77
	assign leaf[1098] = !f[190] && !f[130] && f[406] && f[325]; // c5t775i77
	assign leaf[1099] = !f[190] && f[130] && !f[215] && !f[154]; // c5t775i77
	assign leaf[1100] = !f[190] && f[130] && !f[215] && f[154]; // c5t775i77
	assign leaf[1101] = !f[190] && f[130] && f[215] && !f[239]; // c5t775i77
	assign leaf[1102] = !f[190] && f[130] && f[215] && f[239]; // c5t775i77
	assign leaf[1103] = f[190] && !f[214] && !f[540] && !f[492]; // c5t775i77
	assign leaf[1104] = f[190] && !f[214] && !f[540] && f[492]; // c5t775i77
	assign leaf[1105] = f[190] && !f[214] && f[540] && !f[625]; // c5t775i77
	assign leaf[1106] = f[190] && !f[214] && f[540] && f[625]; // c5t775i77
	assign leaf[1107] = f[190] && f[214] && !f[275] && !f[160]; // c5t775i77
	assign leaf[1108] = f[190] && f[214] && !f[275] && f[160]; // c5t775i77
	assign leaf[1109] = f[190] && f[214] && f[275] && !f[270]; // c5t775i77
	assign leaf[1110] = f[190] && f[214] && f[275] && f[270]; // c5t775i77
	assign leaf[1111] = !f[99] && !f[153] && !f[102] && !f[687]; // c5t785i78
	assign leaf[1112] = !f[99] && !f[153] && !f[102] && f[687]; // c5t785i78
	assign leaf[1113] = !f[99] && !f[153] && f[102] && !f[464]; // c5t785i78
	assign leaf[1114] = !f[99] && !f[153] && f[102] && f[464]; // c5t785i78
	assign leaf[1115] = !f[99] && f[153] && !f[263] && !f[268]; // c5t785i78
	assign leaf[1116] = !f[99] && f[153] && !f[263] && f[268]; // c5t785i78
	assign leaf[1117] = !f[99] && f[153] && f[263] && !f[373]; // c5t785i78
	assign leaf[1118] = !f[99] && f[153] && f[263] && f[373]; // c5t785i78
	assign leaf[1119] = f[99] && !f[181] && !f[294] && !f[289]; // c5t785i78
	assign leaf[1120] = f[99] && !f[181] && !f[294] && f[289]; // c5t785i78
	assign leaf[1121] = f[99] && !f[181] && f[294]; // c5t785i78
	assign leaf[1122] = f[99] && f[181] && !f[458] && !f[237]; // c5t785i78
	assign leaf[1123] = f[99] && f[181] && !f[458] && f[237]; // c5t785i78
	assign leaf[1124] = f[99] && f[181] && f[458]; // c5t785i78
	assign leaf[1125] = !f[411] && !f[468] && !f[354] && !f[301]; // c5t795i79
	assign leaf[1126] = !f[411] && !f[468] && !f[354] && f[301]; // c5t795i79
	assign leaf[1127] = !f[411] && !f[468] && f[354] && !f[324]; // c5t795i79
	assign leaf[1128] = !f[411] && !f[468] && f[354] && f[324]; // c5t795i79
	assign leaf[1129] = !f[411] && f[468] && !f[691] && !f[216]; // c5t795i79
	assign leaf[1130] = !f[411] && f[468] && !f[691] && f[216]; // c5t795i79
	assign leaf[1131] = !f[411] && f[468] && f[691]; // c5t795i79
	assign leaf[1132] = f[411] && !f[523] && !f[149] && !f[374]; // c5t795i79
	assign leaf[1133] = f[411] && !f[523] && !f[149] && f[374]; // c5t795i79
	assign leaf[1134] = f[411] && !f[523] && f[149] && !f[654]; // c5t795i79
	assign leaf[1135] = f[411] && !f[523] && f[149] && f[654]; // c5t795i79
	assign leaf[1136] = f[411] && f[523] && !f[187] && !f[157]; // c5t795i79
	assign leaf[1137] = f[411] && f[523] && !f[187] && f[157]; // c5t795i79
	assign leaf[1138] = f[411] && f[523] && f[187] && !f[237]; // c5t795i79
	assign leaf[1139] = f[411] && f[523] && f[187] && f[237]; // c5t795i79
	assign leaf[1140] = !f[612] && !f[484] && !f[134] && !f[429]; // c5t805i80
	assign leaf[1141] = !f[612] && !f[484] && !f[134] && f[429]; // c5t805i80
	assign leaf[1142] = !f[612] && !f[484] && f[134] && !f[191]; // c5t805i80
	assign leaf[1143] = !f[612] && !f[484] && f[134] && f[191]; // c5t805i80
	assign leaf[1144] = !f[612] && f[484] && !f[429] && !f[459]; // c5t805i80
	assign leaf[1145] = !f[612] && f[484] && !f[429] && f[459]; // c5t805i80
	assign leaf[1146] = !f[612] && f[484] && f[429] && !f[540]; // c5t805i80
	assign leaf[1147] = !f[612] && f[484] && f[429] && f[540]; // c5t805i80
	assign leaf[1148] = f[612]; // c5t805i80
	assign leaf[1149] = !f[411] && !f[440] && !f[357] && !f[325]; // c5t815i81
	assign leaf[1150] = !f[411] && !f[440] && !f[357] && f[325]; // c5t815i81
	assign leaf[1151] = !f[411] && !f[440] && f[357] && !f[272]; // c5t815i81
	assign leaf[1152] = !f[411] && !f[440] && f[357] && f[272]; // c5t815i81
	assign leaf[1153] = !f[411] && f[440] && !f[635] && !f[319]; // c5t815i81
	assign leaf[1154] = !f[411] && f[440] && !f[635] && f[319]; // c5t815i81
	assign leaf[1155] = !f[411] && f[440] && f[635] && !f[210]; // c5t815i81
	assign leaf[1156] = !f[411] && f[440] && f[635] && f[210]; // c5t815i81
	assign leaf[1157] = f[411] && !f[329] && !f[185] && !f[127]; // c5t815i81
	assign leaf[1158] = f[411] && !f[329] && !f[185] && f[127]; // c5t815i81
	assign leaf[1159] = f[411] && !f[329] && f[185] && !f[271]; // c5t815i81
	assign leaf[1160] = f[411] && !f[329] && f[185] && f[271]; // c5t815i81
	assign leaf[1161] = f[411] && f[329] && !f[552]; // c5t815i81
	assign leaf[1162] = f[411] && f[329] && f[552]; // c5t815i81
	assign leaf[1163] = !f[402] && !f[187] && !f[239] && !f[128]; // c5t825i82
	assign leaf[1164] = !f[402] && !f[187] && !f[239] && f[128]; // c5t825i82
	assign leaf[1165] = !f[402] && !f[187] && f[239] && !f[244]; // c5t825i82
	assign leaf[1166] = !f[402] && !f[187] && f[239] && f[244]; // c5t825i82
	assign leaf[1167] = !f[402] && f[187] && !f[211] && !f[215]; // c5t825i82
	assign leaf[1168] = !f[402] && f[187] && !f[211] && f[215]; // c5t825i82
	assign leaf[1169] = !f[402] && f[187] && f[211] && !f[299]; // c5t825i82
	assign leaf[1170] = !f[402] && f[187] && f[211] && f[299]; // c5t825i82
	assign leaf[1171] = f[402] && !f[484] && !f[568] && !f[491]; // c5t825i82
	assign leaf[1172] = f[402] && !f[484] && !f[568] && f[491]; // c5t825i82
	assign leaf[1173] = f[402] && !f[484] && f[568] && !f[319]; // c5t825i82
	assign leaf[1174] = f[402] && !f[484] && f[568] && f[319]; // c5t825i82
	assign leaf[1175] = f[402] && f[484] && !f[625] && !f[638]; // c5t825i82
	assign leaf[1176] = f[402] && f[484] && !f[625] && f[638]; // c5t825i82
	assign leaf[1177] = f[402] && f[484] && f[625] && !f[467]; // c5t825i82
	assign leaf[1178] = f[402] && f[484] && f[625] && f[467]; // c5t825i82
	assign leaf[1179] = !f[276] && !f[380] && !f[681] && !f[521]; // c5t835i83
	assign leaf[1180] = !f[276] && !f[380] && !f[681] && f[521]; // c5t835i83
	assign leaf[1181] = !f[276] && !f[380] && f[681] && !f[548]; // c5t835i83
	assign leaf[1182] = !f[276] && !f[380] && f[681] && f[548]; // c5t835i83
	assign leaf[1183] = !f[276] && f[380] && !f[328] && !f[131]; // c5t835i83
	assign leaf[1184] = !f[276] && f[380] && !f[328] && f[131]; // c5t835i83
	assign leaf[1185] = !f[276] && f[380] && f[328] && !f[407]; // c5t835i83
	assign leaf[1186] = !f[276] && f[380] && f[328] && f[407]; // c5t835i83
	assign leaf[1187] = f[276] && !f[273]; // c5t835i83
	assign leaf[1188] = f[276] && f[273] && !f[234] && !f[351]; // c5t835i83
	assign leaf[1189] = f[276] && f[273] && !f[234] && f[351]; // c5t835i83
	assign leaf[1190] = f[276] && f[273] && f[234]; // c5t835i83
	assign leaf[1191] = !f[216] && !f[322] && !f[599] && !f[524]; // c5t845i84
	assign leaf[1192] = !f[216] && !f[322] && !f[599] && f[524]; // c5t845i84
	assign leaf[1193] = !f[216] && !f[322] && f[599] && !f[242]; // c5t845i84
	assign leaf[1194] = !f[216] && !f[322] && f[599] && f[242]; // c5t845i84
	assign leaf[1195] = !f[216] && f[322] && !f[267] && !f[242]; // c5t845i84
	assign leaf[1196] = !f[216] && f[322] && !f[267] && f[242]; // c5t845i84
	assign leaf[1197] = !f[216] && f[322] && f[267] && !f[299]; // c5t845i84
	assign leaf[1198] = !f[216] && f[322] && f[267] && f[299]; // c5t845i84
	assign leaf[1199] = f[216] && !f[299] && !f[370] && !f[213]; // c5t845i84
	assign leaf[1200] = f[216] && !f[299] && !f[370] && f[213]; // c5t845i84
	assign leaf[1201] = f[216] && !f[299] && f[370] && !f[662]; // c5t845i84
	assign leaf[1202] = f[216] && !f[299] && f[370] && f[662]; // c5t845i84
	assign leaf[1203] = f[216] && f[299] && !f[268]; // c5t845i84
	assign leaf[1204] = f[216] && f[299] && f[268] && !f[272]; // c5t845i84
	assign leaf[1205] = f[216] && f[299] && f[268] && f[272]; // c5t845i84
	assign leaf[1206] = !f[717] && !f[577] && !f[432] && !f[411]; // c5t855i85
	assign leaf[1207] = !f[717] && !f[577] && !f[432] && f[411]; // c5t855i85
	assign leaf[1208] = !f[717] && !f[577] && f[432] && !f[330]; // c5t855i85
	assign leaf[1209] = !f[717] && !f[577] && f[432] && f[330]; // c5t855i85
	assign leaf[1210] = !f[717] && f[577] && !f[397] && !f[216]; // c5t855i85
	assign leaf[1211] = !f[717] && f[577] && !f[397] && f[216]; // c5t855i85
	assign leaf[1212] = !f[717] && f[577] && f[397] && !f[353]; // c5t855i85
	assign leaf[1213] = !f[717] && f[577] && f[397] && f[353]; // c5t855i85
	assign leaf[1214] = f[717] && !f[351] && !f[577]; // c5t855i85
	assign leaf[1215] = f[717] && !f[351] && f[577]; // c5t855i85
	assign leaf[1216] = f[717] && f[351]; // c5t855i85
	assign leaf[1217] = !f[685] && !f[521] && !f[205] && !f[318]; // c5t865i86
	assign leaf[1218] = !f[685] && !f[521] && !f[205] && f[318]; // c5t865i86
	assign leaf[1219] = !f[685] && !f[521] && f[205] && !f[375]; // c5t865i86
	assign leaf[1220] = !f[685] && !f[521] && f[205] && f[375]; // c5t865i86
	assign leaf[1221] = !f[685] && f[521] && !f[234] && !f[548]; // c5t865i86
	assign leaf[1222] = !f[685] && f[521] && !f[234] && f[548]; // c5t865i86
	assign leaf[1223] = !f[685] && f[521] && f[234] && !f[127]; // c5t865i86
	assign leaf[1224] = !f[685] && f[521] && f[234] && f[127]; // c5t865i86
	assign leaf[1225] = f[685] && !f[546] && !f[290] && !f[294]; // c5t865i86
	assign leaf[1226] = f[685] && !f[546] && !f[290] && f[294]; // c5t865i86
	assign leaf[1227] = f[685] && !f[546] && f[290] && !f[174]; // c5t865i86
	assign leaf[1228] = f[685] && !f[546] && f[290] && f[174]; // c5t865i86
	assign leaf[1229] = f[685] && f[546] && !f[210]; // c5t865i86
	assign leaf[1230] = f[685] && f[546] && f[210] && !f[274]; // c5t865i86
	assign leaf[1231] = f[685] && f[546] && f[210] && f[274]; // c5t865i86
	assign leaf[1232] = !f[333] && !f[622] && !f[598] && !f[654]; // c5t875i87
	assign leaf[1233] = !f[333] && !f[622] && !f[598] && f[654]; // c5t875i87
	assign leaf[1234] = !f[333] && !f[622] && f[598] && !f[397]; // c5t875i87
	assign leaf[1235] = !f[333] && !f[622] && f[598] && f[397]; // c5t875i87
	assign leaf[1236] = !f[333] && f[622] && !f[540] && !f[179]; // c5t875i87
	assign leaf[1237] = !f[333] && f[622] && !f[540] && f[179]; // c5t875i87
	assign leaf[1238] = !f[333] && f[622] && f[540] && !f[537]; // c5t875i87
	assign leaf[1239] = !f[333] && f[622] && f[540] && f[537]; // c5t875i87
	assign leaf[1240] = f[333]; // c5t875i87
	assign leaf[1241] = !f[492] && !f[490] && !f[510] && !f[99]; // c5t885i88
	assign leaf[1242] = !f[492] && !f[490] && !f[510] && f[99]; // c5t885i88
	assign leaf[1243] = !f[492] && !f[490] && f[510] && !f[625]; // c5t885i88
	assign leaf[1244] = !f[492] && !f[490] && f[510] && f[625]; // c5t885i88
	assign leaf[1245] = !f[492] && f[490] && !f[261] && !f[331]; // c5t885i88
	assign leaf[1246] = !f[492] && f[490] && !f[261] && f[331]; // c5t885i88
	assign leaf[1247] = !f[492] && f[490] && f[261] && !f[319]; // c5t885i88
	assign leaf[1248] = !f[492] && f[490] && f[261] && f[319]; // c5t885i88
	assign leaf[1249] = f[492] && !f[625] && !f[511] && !f[684]; // c5t885i88
	assign leaf[1250] = f[492] && !f[625] && !f[511] && f[684]; // c5t885i88
	assign leaf[1251] = f[492] && !f[625] && f[511] && !f[538]; // c5t885i88
	assign leaf[1252] = f[492] && !f[625] && f[511] && f[538]; // c5t885i88
	assign leaf[1253] = f[492] && f[625] && !f[321] && !f[409]; // c5t885i88
	assign leaf[1254] = f[492] && f[625] && !f[321] && f[409]; // c5t885i88
	assign leaf[1255] = f[492] && f[625] && f[321] && !f[296]; // c5t885i88
	assign leaf[1256] = f[492] && f[625] && f[321] && f[296]; // c5t885i88
	assign leaf[1257] = !f[351] && !f[454] && !f[296] && !f[327]; // c5t895i89
	assign leaf[1258] = !f[351] && !f[454] && !f[296] && f[327]; // c5t895i89
	assign leaf[1259] = !f[351] && !f[454] && f[296] && !f[184]; // c5t895i89
	assign leaf[1260] = !f[351] && !f[454] && f[296] && f[184]; // c5t895i89
	assign leaf[1261] = !f[351] && f[454] && !f[457] && !f[427]; // c5t895i89
	assign leaf[1262] = !f[351] && f[454] && !f[457] && f[427]; // c5t895i89
	assign leaf[1263] = !f[351] && f[454] && f[457] && !f[374]; // c5t895i89
	assign leaf[1264] = !f[351] && f[454] && f[457] && f[374]; // c5t895i89
	assign leaf[1265] = f[351] && !f[406] && !f[155] && !f[552]; // c5t895i89
	assign leaf[1266] = f[351] && !f[406] && !f[155] && f[552]; // c5t895i89
	assign leaf[1267] = f[351] && !f[406] && f[155] && !f[240]; // c5t895i89
	assign leaf[1268] = f[351] && !f[406] && f[155] && f[240]; // c5t895i89
	assign leaf[1269] = f[351] && f[406] && !f[540] && !f[348]; // c5t895i89
	assign leaf[1270] = f[351] && f[406] && !f[540] && f[348]; // c5t895i89
	assign leaf[1271] = f[351] && f[406] && f[540] && !f[325]; // c5t895i89
	assign leaf[1272] = f[351] && f[406] && f[540] && f[325]; // c5t895i89
	assign leaf[1273] = !f[119] && !f[322] && !f[519] && !f[517]; // c5t905i90
	assign leaf[1274] = !f[119] && !f[322] && !f[519] && f[517]; // c5t905i90
	assign leaf[1275] = !f[119] && !f[322] && f[519] && !f[295]; // c5t905i90
	assign leaf[1276] = !f[119] && !f[322] && f[519] && f[295]; // c5t905i90
	assign leaf[1277] = !f[119] && f[322] && !f[491] && !f[462]; // c5t905i90
	assign leaf[1278] = !f[119] && f[322] && !f[491] && f[462]; // c5t905i90
	assign leaf[1279] = !f[119] && f[322] && f[491] && !f[265]; // c5t905i90
	assign leaf[1280] = !f[119] && f[322] && f[491] && f[265]; // c5t905i90
	assign leaf[1281] = f[119] && !f[609]; // c5t905i90
	assign leaf[1282] = f[119] && f[609]; // c5t905i90
	assign leaf[1283] = !f[485] && !f[291] && !f[596] && !f[266]; // c5t915i91
	assign leaf[1284] = !f[485] && !f[291] && !f[596] && f[266]; // c5t915i91
	assign leaf[1285] = !f[485] && !f[291] && f[596] && !f[235]; // c5t915i91
	assign leaf[1286] = !f[485] && !f[291] && f[596] && f[235]; // c5t915i91
	assign leaf[1287] = !f[485] && f[291] && !f[207] && !f[407]; // c5t915i91
	assign leaf[1288] = !f[485] && f[291] && !f[207] && f[407]; // c5t915i91
	assign leaf[1289] = !f[485] && f[291] && f[207] && !f[235]; // c5t915i91
	assign leaf[1290] = !f[485] && f[291] && f[207] && f[235]; // c5t915i91
	assign leaf[1291] = f[485] && !f[407] && !f[136] && !f[541]; // c5t915i91
	assign leaf[1292] = f[485] && !f[407] && !f[136] && f[541]; // c5t915i91
	assign leaf[1293] = f[485] && !f[407] && f[136]; // c5t915i91
	assign leaf[1294] = f[485] && f[407] && !f[515] && !f[569]; // c5t915i91
	assign leaf[1295] = f[485] && f[407] && !f[515] && f[569]; // c5t915i91
	assign leaf[1296] = f[485] && f[407] && f[515] && !f[577]; // c5t915i91
	assign leaf[1297] = f[485] && f[407] && f[515] && f[577]; // c5t915i91
	assign leaf[1298] = !f[627] && !f[428] && !f[271] && !f[184]; // c5t925i92
	assign leaf[1299] = !f[627] && !f[428] && !f[271] && f[184]; // c5t925i92
	assign leaf[1300] = !f[627] && !f[428] && f[271] && !f[269]; // c5t925i92
	assign leaf[1301] = !f[627] && !f[428] && f[271] && f[269]; // c5t925i92
	assign leaf[1302] = !f[627] && f[428] && !f[290] && !f[510]; // c5t925i92
	assign leaf[1303] = !f[627] && f[428] && !f[290] && f[510]; // c5t925i92
	assign leaf[1304] = !f[627] && f[428] && f[290] && !f[128]; // c5t925i92
	assign leaf[1305] = !f[627] && f[428] && f[290] && f[128]; // c5t925i92
	assign leaf[1306] = f[627] && !f[463] && !f[234] && !f[290]; // c5t925i92
	assign leaf[1307] = f[627] && !f[463] && !f[234] && f[290]; // c5t925i92
	assign leaf[1308] = f[627] && !f[463] && f[234] && !f[269]; // c5t925i92
	assign leaf[1309] = f[627] && !f[463] && f[234] && f[269]; // c5t925i92
	assign leaf[1310] = f[627] && f[463] && !f[547] && !f[321]; // c5t925i92
	assign leaf[1311] = f[627] && f[463] && !f[547] && f[321]; // c5t925i92
	assign leaf[1312] = f[627] && f[463] && f[547] && !f[384]; // c5t925i92
	assign leaf[1313] = f[627] && f[463] && f[547] && f[384]; // c5t925i92
	assign leaf[1314] = !f[276] && !f[434] && !f[520] && !f[322]; // c5t935i93
	assign leaf[1315] = !f[276] && !f[434] && !f[520] && f[322]; // c5t935i93
	assign leaf[1316] = !f[276] && !f[434] && f[520] && !f[264]; // c5t935i93
	assign leaf[1317] = !f[276] && !f[434] && f[520] && f[264]; // c5t935i93
	assign leaf[1318] = !f[276] && f[434] && !f[325] && !f[215]; // c5t935i93
	assign leaf[1319] = !f[276] && f[434] && !f[325] && f[215]; // c5t935i93
	assign leaf[1320] = !f[276] && f[434] && f[325] && !f[352]; // c5t935i93
	assign leaf[1321] = !f[276] && f[434] && f[325] && f[352]; // c5t935i93
	assign leaf[1322] = f[276] && !f[273]; // c5t935i93
	assign leaf[1323] = f[276] && f[273] && !f[262] && !f[351]; // c5t935i93
	assign leaf[1324] = f[276] && f[273] && !f[262] && f[351]; // c5t935i93
	assign leaf[1325] = f[276] && f[273] && f[262]; // c5t935i93
	assign leaf[1326] = !f[612] && !f[147] && !f[258] && !f[155]; // c5t945i94
	assign leaf[1327] = !f[612] && !f[147] && !f[258] && f[155]; // c5t945i94
	assign leaf[1328] = !f[612] && !f[147] && f[258] && !f[399]; // c5t945i94
	assign leaf[1329] = !f[612] && !f[147] && f[258] && f[399]; // c5t945i94
	assign leaf[1330] = !f[612] && f[147] && !f[204] && !f[208]; // c5t945i94
	assign leaf[1331] = !f[612] && f[147] && !f[204] && f[208]; // c5t945i94
	assign leaf[1332] = !f[612] && f[147] && f[204] && !f[498]; // c5t945i94
	assign leaf[1333] = !f[612] && f[147] && f[204] && f[498]; // c5t945i94
	assign leaf[1334] = f[612]; // c5t945i94
	assign leaf[1335] = !f[636] && !f[177] && !f[315] && !f[232]; // c5t955i95
	assign leaf[1336] = !f[636] && !f[177] && !f[315] && f[232]; // c5t955i95
	assign leaf[1337] = !f[636] && !f[177] && f[315] && !f[204]; // c5t955i95
	assign leaf[1338] = !f[636] && !f[177] && f[315] && f[204]; // c5t955i95
	assign leaf[1339] = !f[636] && f[177] && !f[128] && !f[206]; // c5t955i95
	assign leaf[1340] = !f[636] && f[177] && !f[128] && f[206]; // c5t955i95
	assign leaf[1341] = !f[636] && f[177] && f[128] && !f[261]; // c5t955i95
	assign leaf[1342] = !f[636] && f[177] && f[128] && f[261]; // c5t955i95
	assign leaf[1343] = f[636] && !f[344] && !f[406] && !f[266]; // c5t955i95
	assign leaf[1344] = f[636] && !f[344] && !f[406] && f[266]; // c5t955i95
	assign leaf[1345] = f[636] && !f[344] && f[406] && !f[598]; // c5t955i95
	assign leaf[1346] = f[636] && !f[344] && f[406] && f[598]; // c5t955i95
	assign leaf[1347] = f[636] && f[344] && !f[260] && !f[378]; // c5t955i95
	assign leaf[1348] = f[636] && f[344] && !f[260] && f[378]; // c5t955i95
	assign leaf[1349] = f[636] && f[344] && f[260] && !f[660]; // c5t955i95
	assign leaf[1350] = f[636] && f[344] && f[260] && f[660]; // c5t955i95
	assign leaf[1351] = !f[380] && !f[686] && !f[549] && !f[293]; // c5t965i96
	assign leaf[1352] = !f[380] && !f[686] && !f[549] && f[293]; // c5t965i96
	assign leaf[1353] = !f[380] && !f[686] && f[549] && !f[427]; // c5t965i96
	assign leaf[1354] = !f[380] && !f[686] && f[549] && f[427]; // c5t965i96
	assign leaf[1355] = !f[380] && f[686] && !f[289] && !f[296]; // c5t965i96
	assign leaf[1356] = !f[380] && f[686] && !f[289] && f[296]; // c5t965i96
	assign leaf[1357] = !f[380] && f[686] && f[289] && !f[572]; // c5t965i96
	assign leaf[1358] = !f[380] && f[686] && f[289] && f[572]; // c5t965i96
	assign leaf[1359] = f[380] && !f[248] && !f[342] && !f[522]; // c5t965i96
	assign leaf[1360] = f[380] && !f[248] && !f[342] && f[522]; // c5t965i96
	assign leaf[1361] = f[380] && !f[248] && f[342] && !f[347]; // c5t965i96
	assign leaf[1362] = f[380] && !f[248] && f[342] && f[347]; // c5t965i96
	assign leaf[1363] = f[380] && f[248] && !f[219]; // c5t965i96
	assign leaf[1364] = f[380] && f[248] && f[219]; // c5t965i96
	assign leaf[1365] = !f[707] && !f[424] && !f[508] && !f[322]; // c5t975i97
	assign leaf[1366] = !f[707] && !f[424] && !f[508] && f[322]; // c5t975i97
	assign leaf[1367] = !f[707] && !f[424] && f[508] && !f[301]; // c5t975i97
	assign leaf[1368] = !f[707] && !f[424] && f[508] && f[301]; // c5t975i97
	assign leaf[1369] = !f[707] && f[424] && !f[357]; // c5t975i97
	assign leaf[1370] = !f[707] && f[424] && f[357]; // c5t975i97
	assign leaf[1371] = f[707]; // c5t975i97
	assign leaf[1372] = !f[411] && !f[158] && !f[434] && !f[270]; // c5t985i98
	assign leaf[1373] = !f[411] && !f[158] && !f[434] && f[270]; // c5t985i98
	assign leaf[1374] = !f[411] && !f[158] && f[434] && !f[352]; // c5t985i98
	assign leaf[1375] = !f[411] && !f[158] && f[434] && f[352]; // c5t985i98
	assign leaf[1376] = !f[411] && f[158] && !f[243] && !f[245]; // c5t985i98
	assign leaf[1377] = !f[411] && f[158] && !f[243] && f[245]; // c5t985i98
	assign leaf[1378] = !f[411] && f[158] && f[243] && !f[434]; // c5t985i98
	assign leaf[1379] = !f[411] && f[158] && f[243] && f[434]; // c5t985i98
	assign leaf[1380] = f[411] && !f[300] && !f[593] && !f[131]; // c5t985i98
	assign leaf[1381] = f[411] && !f[300] && !f[593] && f[131]; // c5t985i98
	assign leaf[1382] = f[411] && !f[300] && f[593] && !f[237]; // c5t985i98
	assign leaf[1383] = f[411] && !f[300] && f[593] && f[237]; // c5t985i98
	assign leaf[1384] = f[411] && f[300] && !f[383]; // c5t985i98
	assign leaf[1385] = f[411] && f[300] && f[383] && !f[356]; // c5t985i98
	assign leaf[1386] = f[411] && f[300] && f[383] && f[356]; // c5t985i98
	assign leaf[1387] = !f[297] && !f[215] && !f[266] && !f[127]; // c5t995i99
	assign leaf[1388] = !f[297] && !f[215] && !f[266] && f[127]; // c5t995i99
	assign leaf[1389] = !f[297] && !f[215] && f[266] && !f[623]; // c5t995i99
	assign leaf[1390] = !f[297] && !f[215] && f[266] && f[623]; // c5t995i99
	assign leaf[1391] = !f[297] && f[215] && !f[372] && !f[299]; // c5t995i99
	assign leaf[1392] = !f[297] && f[215] && !f[372] && f[299]; // c5t995i99
	assign leaf[1393] = !f[297] && f[215] && f[372] && !f[454]; // c5t995i99
	assign leaf[1394] = !f[297] && f[215] && f[372] && f[454]; // c5t995i99
	assign leaf[1395] = f[297] && !f[295] && !f[414] && !f[267]; // c5t995i99
	assign leaf[1396] = f[297] && !f[295] && !f[414] && f[267]; // c5t995i99
	assign leaf[1397] = f[297] && !f[295] && f[414]; // c5t995i99
	assign leaf[1398] = f[297] && f[295] && !f[242] && !f[342]; // c5t995i99
	assign leaf[1399] = f[297] && f[295] && !f[242] && f[342]; // c5t995i99
	assign leaf[1400] = f[297] && f[295] && f[242] && !f[156]; // c5t995i99
	assign leaf[1401] = f[297] && f[295] && f[242] && f[156]; // c5t995i99
endmodule

module decision_tree_leaves_6(input logic [0:783] f, output logic [0:1336] leaf);
	assign leaf[0] = !f[101] && !f[98] && !f[103] && !f[95]; // c6t6i0
	assign leaf[1] = !f[101] && !f[98] && !f[103] && f[95]; // c6t6i0
	assign leaf[2] = !f[101] && !f[98] && f[103] && !f[244]; // c6t6i0
	assign leaf[3] = !f[101] && !f[98] && f[103] && f[244]; // c6t6i0
	assign leaf[4] = !f[101] && f[98] && !f[213] && !f[267]; // c6t6i0
	assign leaf[5] = !f[101] && f[98] && !f[213] && f[267]; // c6t6i0
	assign leaf[6] = !f[101] && f[98] && f[213] && !f[291]; // c6t6i0
	assign leaf[7] = !f[101] && f[98] && f[213] && f[291]; // c6t6i0
	assign leaf[8] = f[101] && !f[243] && !f[594] && !f[269]; // c6t6i0
	assign leaf[9] = f[101] && !f[243] && !f[594] && f[269]; // c6t6i0
	assign leaf[10] = f[101] && !f[243] && f[594] && !f[292]; // c6t6i0
	assign leaf[11] = f[101] && !f[243] && f[594] && f[292]; // c6t6i0
	assign leaf[12] = f[101] && f[243] && !f[317] && !f[318]; // c6t6i0
	assign leaf[13] = f[101] && f[243] && !f[317] && f[318]; // c6t6i0
	assign leaf[14] = f[101] && f[243] && f[317] && !f[461]; // c6t6i0
	assign leaf[15] = f[101] && f[243] && f[317] && f[461]; // c6t6i0
	assign leaf[16] = !f[514] && !f[101] && !f[70] && !f[105]; // c6t16i1
	assign leaf[17] = !f[514] && !f[101] && !f[70] && f[105]; // c6t16i1
	assign leaf[18] = !f[514] && !f[101] && f[70] && !f[156]; // c6t16i1
	assign leaf[19] = !f[514] && !f[101] && f[70] && f[156]; // c6t16i1
	assign leaf[20] = !f[514] && f[101] && !f[625] && !f[237]; // c6t16i1
	assign leaf[21] = !f[514] && f[101] && !f[625] && f[237]; // c6t16i1
	assign leaf[22] = !f[514] && f[101] && f[625] && !f[414]; // c6t16i1
	assign leaf[23] = !f[514] && f[101] && f[625] && f[414]; // c6t16i1
	assign leaf[24] = f[514] && !f[242] && !f[245] && !f[268]; // c6t16i1
	assign leaf[25] = f[514] && !f[242] && !f[245] && f[268]; // c6t16i1
	assign leaf[26] = f[514] && !f[242] && f[245] && !f[120]; // c6t16i1
	assign leaf[27] = f[514] && !f[242] && f[245] && f[120]; // c6t16i1
	assign leaf[28] = f[514] && f[242] && !f[105] && !f[135]; // c6t16i1
	assign leaf[29] = f[514] && f[242] && !f[105] && f[135]; // c6t16i1
	assign leaf[30] = f[514] && f[242] && f[105] && !f[325]; // c6t16i1
	assign leaf[31] = f[514] && f[242] && f[105] && f[325]; // c6t16i1
	assign leaf[32] = !f[543] && !f[104] && !f[101] && !f[69]; // c6t26i2
	assign leaf[33] = !f[543] && !f[104] && !f[101] && f[69]; // c6t26i2
	assign leaf[34] = !f[543] && !f[104] && f[101] && !f[402]; // c6t26i2
	assign leaf[35] = !f[543] && !f[104] && f[101] && f[402]; // c6t26i2
	assign leaf[36] = !f[543] && f[104] && !f[541] && !f[266]; // c6t26i2
	assign leaf[37] = !f[543] && f[104] && !f[541] && f[266]; // c6t26i2
	assign leaf[38] = !f[543] && f[104] && f[541] && !f[103]; // c6t26i2
	assign leaf[39] = !f[543] && f[104] && f[541] && f[103]; // c6t26i2
	assign leaf[40] = f[543] && !f[242] && !f[655] && !f[216]; // c6t26i2
	assign leaf[41] = f[543] && !f[242] && !f[655] && f[216]; // c6t26i2
	assign leaf[42] = f[543] && !f[242] && f[655] && !f[131]; // c6t26i2
	assign leaf[43] = f[543] && !f[242] && f[655] && f[131]; // c6t26i2
	assign leaf[44] = f[543] && f[242] && !f[106] && !f[104]; // c6t26i2
	assign leaf[45] = f[543] && f[242] && !f[106] && f[104]; // c6t26i2
	assign leaf[46] = f[543] && f[242] && f[106] && !f[325]; // c6t26i2
	assign leaf[47] = f[543] && f[242] && f[106] && f[325]; // c6t26i2
	assign leaf[48] = !f[543] && !f[570] && !f[68] && !f[70]; // c6t36i3
	assign leaf[49] = !f[543] && !f[570] && !f[68] && f[70]; // c6t36i3
	assign leaf[50] = !f[543] && !f[570] && f[68]; // c6t36i3
	assign leaf[51] = !f[543] && f[570] && !f[271] && !f[457]; // c6t36i3
	assign leaf[52] = !f[543] && f[570] && !f[271] && f[457]; // c6t36i3
	assign leaf[53] = !f[543] && f[570] && f[271] && !f[92]; // c6t36i3
	assign leaf[54] = !f[543] && f[570] && f[271] && f[92]; // c6t36i3
	assign leaf[55] = f[543] && !f[242] && !f[575] && !f[296]; // c6t36i3
	assign leaf[56] = f[543] && !f[242] && !f[575] && f[296]; // c6t36i3
	assign leaf[57] = f[543] && !f[242] && f[575] && !f[625]; // c6t36i3
	assign leaf[58] = f[543] && !f[242] && f[575] && f[625]; // c6t36i3
	assign leaf[59] = f[543] && f[242] && !f[105] && !f[457]; // c6t36i3
	assign leaf[60] = f[543] && f[242] && !f[105] && f[457]; // c6t36i3
	assign leaf[61] = f[543] && f[242] && f[105] && !f[298]; // c6t36i3
	assign leaf[62] = f[543] && f[242] && f[105] && f[298]; // c6t36i3
	assign leaf[63] = !f[514] && !f[512] && !f[515] && !f[387]; // c6t46i4
	assign leaf[64] = !f[514] && !f[512] && !f[515] && f[387]; // c6t46i4
	assign leaf[65] = !f[514] && !f[512] && f[515] && !f[431]; // c6t46i4
	assign leaf[66] = !f[514] && !f[512] && f[515] && f[431]; // c6t46i4
	assign leaf[67] = !f[514] && f[512] && !f[243] && !f[269]; // c6t46i4
	assign leaf[68] = !f[514] && f[512] && !f[243] && f[269]; // c6t46i4
	assign leaf[69] = !f[514] && f[512] && f[243] && !f[135]; // c6t46i4
	assign leaf[70] = !f[514] && f[512] && f[243] && f[135]; // c6t46i4
	assign leaf[71] = f[514] && !f[270] && !f[272] && !f[296]; // c6t46i4
	assign leaf[72] = f[514] && !f[270] && !f[272] && f[296]; // c6t46i4
	assign leaf[73] = f[514] && !f[270] && f[272] && !f[388]; // c6t46i4
	assign leaf[74] = f[514] && !f[270] && f[272] && f[388]; // c6t46i4
	assign leaf[75] = f[514] && f[270] && !f[386] && !f[106]; // c6t46i4
	assign leaf[76] = f[514] && f[270] && !f[386] && f[106]; // c6t46i4
	assign leaf[77] = f[514] && f[270] && f[386] && !f[241]; // c6t46i4
	assign leaf[78] = f[514] && f[270] && f[386] && f[241]; // c6t46i4
	assign leaf[79] = !f[270] && !f[543] && !f[541] && !f[516]; // c6t56i5
	assign leaf[80] = !f[270] && !f[543] && !f[541] && f[516]; // c6t56i5
	assign leaf[81] = !f[270] && !f[543] && f[541] && !f[244]; // c6t56i5
	assign leaf[82] = !f[270] && !f[543] && f[541] && f[244]; // c6t56i5
	assign leaf[83] = !f[270] && f[543] && !f[574] && !f[601]; // c6t56i5
	assign leaf[84] = !f[270] && f[543] && !f[574] && f[601]; // c6t56i5
	assign leaf[85] = !f[270] && f[543] && f[574] && !f[245]; // c6t56i5
	assign leaf[86] = !f[270] && f[543] && f[574] && f[245]; // c6t56i5
	assign leaf[87] = f[270] && !f[92] && !f[136] && !f[94]; // c6t56i5
	assign leaf[88] = f[270] && !f[92] && !f[136] && f[94]; // c6t56i5
	assign leaf[89] = f[270] && !f[92] && f[136] && !f[429]; // c6t56i5
	assign leaf[90] = f[270] && !f[92] && f[136] && f[429]; // c6t56i5
	assign leaf[91] = f[270] && f[92] && !f[123] && !f[150]; // c6t56i5
	assign leaf[92] = f[270] && f[92] && !f[123] && f[150]; // c6t56i5
	assign leaf[93] = f[270] && f[92] && f[123]; // c6t56i5
	assign leaf[94] = !f[270] && !f[486] && !f[484] && !f[487]; // c6t66i6
	assign leaf[95] = !f[270] && !f[486] && !f[484] && f[487]; // c6t66i6
	assign leaf[96] = !f[270] && !f[486] && f[484] && !f[244]; // c6t66i6
	assign leaf[97] = !f[270] && !f[486] && f[484] && f[244]; // c6t66i6
	assign leaf[98] = !f[270] && f[486] && !f[272] && !f[296]; // c6t66i6
	assign leaf[99] = !f[270] && f[486] && !f[272] && f[296]; // c6t66i6
	assign leaf[100] = !f[270] && f[486] && f[272] && !f[359]; // c6t66i6
	assign leaf[101] = !f[270] && f[486] && f[272] && f[359]; // c6t66i6
	assign leaf[102] = f[270] && !f[386] && !f[107] && !f[359]; // c6t66i6
	assign leaf[103] = f[270] && !f[386] && !f[107] && f[359]; // c6t66i6
	assign leaf[104] = f[270] && !f[386] && f[107]; // c6t66i6
	assign leaf[105] = f[270] && f[386] && !f[122] && !f[119]; // c6t66i6
	assign leaf[106] = f[270] && f[386] && !f[122] && f[119]; // c6t66i6
	assign leaf[107] = f[270] && f[386] && f[122] && !f[212]; // c6t66i6
	assign leaf[108] = f[270] && f[386] && f[122] && f[212]; // c6t66i6
	assign leaf[109] = !f[242] && !f[572] && !f[388] && !f[131]; // c6t76i7
	assign leaf[110] = !f[242] && !f[572] && !f[388] && f[131]; // c6t76i7
	assign leaf[111] = !f[242] && !f[572] && f[388] && !f[329]; // c6t76i7
	assign leaf[112] = !f[242] && !f[572] && f[388] && f[329]; // c6t76i7
	assign leaf[113] = !f[242] && f[572] && !f[655] && !f[295]; // c6t76i7
	assign leaf[114] = !f[242] && f[572] && !f[655] && f[295]; // c6t76i7
	assign leaf[115] = !f[242] && f[572] && f[655] && !f[131]; // c6t76i7
	assign leaf[116] = !f[242] && f[572] && f[655] && f[131]; // c6t76i7
	assign leaf[117] = f[242] && !f[133] && !f[93] && !f[103]; // c6t76i7
	assign leaf[118] = f[242] && !f[133] && !f[93] && f[103]; // c6t76i7
	assign leaf[119] = f[242] && !f[133] && f[93] && !f[125]; // c6t76i7
	assign leaf[120] = f[242] && !f[133] && f[93] && f[125]; // c6t76i7
	assign leaf[121] = f[242] && f[133] && !f[298] && !f[513]; // c6t76i7
	assign leaf[122] = f[242] && f[133] && !f[298] && f[513]; // c6t76i7
	assign leaf[123] = f[242] && f[133] && f[298] && !f[326]; // c6t76i7
	assign leaf[124] = f[242] && f[133] && f[298] && f[326]; // c6t76i7
	assign leaf[125] = !f[486] && !f[484] && !f[388] && !f[487]; // c6t86i8
	assign leaf[126] = !f[486] && !f[484] && !f[388] && f[487]; // c6t86i8
	assign leaf[127] = !f[486] && !f[484] && f[388] && !f[266]; // c6t86i8
	assign leaf[128] = !f[486] && !f[484] && f[388] && f[266]; // c6t86i8
	assign leaf[129] = !f[486] && f[484] && !f[243] && !f[217]; // c6t86i8
	assign leaf[130] = !f[486] && f[484] && !f[243] && f[217]; // c6t86i8
	assign leaf[131] = !f[486] && f[484] && f[243] && !f[93]; // c6t86i8
	assign leaf[132] = !f[486] && f[484] && f[243] && f[93]; // c6t86i8
	assign leaf[133] = f[486] && !f[271] && !f[402] && !f[414]; // c6t86i8
	assign leaf[134] = f[486] && !f[271] && !f[402] && f[414]; // c6t86i8
	assign leaf[135] = f[486] && !f[271] && f[402] && !f[274]; // c6t86i8
	assign leaf[136] = f[486] && !f[271] && f[402] && f[274]; // c6t86i8
	assign leaf[137] = f[486] && f[271] && !f[121] && !f[96]; // c6t86i8
	assign leaf[138] = f[486] && f[271] && !f[121] && f[96]; // c6t86i8
	assign leaf[139] = f[486] && f[271] && f[121] && !f[185]; // c6t86i8
	assign leaf[140] = f[486] && f[271] && f[121] && f[185]; // c6t86i8
	assign leaf[141] = !f[269] && !f[244] && !f[323] && !f[246]; // c6t96i9
	assign leaf[142] = !f[269] && !f[244] && !f[323] && f[246]; // c6t96i9
	assign leaf[143] = !f[269] && !f[244] && f[323] && !f[430]; // c6t96i9
	assign leaf[144] = !f[269] && !f[244] && f[323] && f[430]; // c6t96i9
	assign leaf[145] = !f[269] && f[244] && !f[355] && !f[513]; // c6t96i9
	assign leaf[146] = !f[269] && f[244] && !f[355] && f[513]; // c6t96i9
	assign leaf[147] = !f[269] && f[244] && f[355] && !f[414]; // c6t96i9
	assign leaf[148] = !f[269] && f[244] && f[355] && f[414]; // c6t96i9
	assign leaf[149] = f[269] && !f[133] && !f[386] && !f[164]; // c6t96i9
	assign leaf[150] = f[269] && !f[133] && !f[386] && f[164]; // c6t96i9
	assign leaf[151] = f[269] && !f[133] && f[386] && !f[239]; // c6t96i9
	assign leaf[152] = f[269] && !f[133] && f[386] && f[239]; // c6t96i9
	assign leaf[153] = f[269] && f[133] && !f[325] && !f[273]; // c6t96i9
	assign leaf[154] = f[269] && f[133] && !f[325] && f[273]; // c6t96i9
	assign leaf[155] = f[269] && f[133] && f[325] && !f[266]; // c6t96i9
	assign leaf[156] = f[269] && f[133] && f[325] && f[266]; // c6t96i9
	assign leaf[157] = !f[269] && !f[243] && !f[549] && !f[323]; // c6t106i10
	assign leaf[158] = !f[269] && !f[243] && !f[549] && f[323]; // c6t106i10
	assign leaf[159] = !f[269] && !f[243] && f[549] && !f[633]; // c6t106i10
	assign leaf[160] = !f[269] && !f[243] && f[549] && f[633]; // c6t106i10
	assign leaf[161] = !f[269] && f[243] && !f[327] && !f[486]; // c6t106i10
	assign leaf[162] = !f[269] && f[243] && !f[327] && f[486]; // c6t106i10
	assign leaf[163] = !f[269] && f[243] && f[327] && !f[358]; // c6t106i10
	assign leaf[164] = !f[269] && f[243] && f[327] && f[358]; // c6t106i10
	assign leaf[165] = f[269] && !f[133] && !f[94] && !f[103]; // c6t106i10
	assign leaf[166] = f[269] && !f[133] && !f[94] && f[103]; // c6t106i10
	assign leaf[167] = f[269] && !f[133] && f[94] && !f[232]; // c6t106i10
	assign leaf[168] = f[269] && !f[133] && f[94] && f[232]; // c6t106i10
	assign leaf[169] = f[269] && f[133] && !f[299] && !f[349]; // c6t106i10
	assign leaf[170] = f[269] && f[133] && !f[299] && f[349]; // c6t106i10
	assign leaf[171] = f[269] && f[133] && f[299]; // c6t106i10
	assign leaf[172] = !f[573] && !f[600] && !f[387] && !f[68]; // c6t116i11
	assign leaf[173] = !f[573] && !f[600] && !f[387] && f[68]; // c6t116i11
	assign leaf[174] = !f[573] && !f[600] && f[387] && !f[520]; // c6t116i11
	assign leaf[175] = !f[573] && !f[600] && f[387] && f[520]; // c6t116i11
	assign leaf[176] = !f[573] && f[600] && !f[458] && !f[427]; // c6t116i11
	assign leaf[177] = !f[573] && f[600] && !f[458] && f[427]; // c6t116i11
	assign leaf[178] = !f[573] && f[600] && f[458] && !f[297]; // c6t116i11
	assign leaf[179] = !f[573] && f[600] && f[458] && f[297]; // c6t116i11
	assign leaf[180] = f[573] && !f[656] && !f[625] && !f[240]; // c6t116i11
	assign leaf[181] = f[573] && !f[656] && !f[625] && f[240]; // c6t116i11
	assign leaf[182] = f[573] && !f[656] && f[625] && !f[107]; // c6t116i11
	assign leaf[183] = f[573] && !f[656] && f[625] && f[107]; // c6t116i11
	assign leaf[184] = f[573] && f[656] && !f[132] && !f[134]; // c6t116i11
	assign leaf[185] = f[573] && f[656] && !f[132] && f[134]; // c6t116i11
	assign leaf[186] = f[573] && f[656] && f[132] && !f[381]; // c6t116i11
	assign leaf[187] = f[573] && f[656] && f[132] && f[381]; // c6t116i11
	assign leaf[188] = !f[269] && !f[654] && !f[576] && !f[548]; // c6t126i12
	assign leaf[189] = !f[269] && !f[654] && !f[576] && f[548]; // c6t126i12
	assign leaf[190] = !f[269] && !f[654] && f[576] && !f[660]; // c6t126i12
	assign leaf[191] = !f[269] && !f[654] && f[576] && f[660]; // c6t126i12
	assign leaf[192] = !f[269] && f[654] && !f[134] && !f[131]; // c6t126i12
	assign leaf[193] = !f[269] && f[654] && !f[134] && f[131]; // c6t126i12
	assign leaf[194] = !f[269] && f[654] && f[134] && !f[353]; // c6t126i12
	assign leaf[195] = !f[269] && f[654] && f[134] && f[353]; // c6t126i12
	assign leaf[196] = f[269] && !f[163] && !f[357] && !f[132]; // c6t126i12
	assign leaf[197] = f[269] && !f[163] && !f[357] && f[132]; // c6t126i12
	assign leaf[198] = f[269] && !f[163] && f[357] && !f[239]; // c6t126i12
	assign leaf[199] = f[269] && !f[163] && f[357] && f[239]; // c6t126i12
	assign leaf[200] = f[269] && f[163] && !f[349]; // c6t126i12
	assign leaf[201] = f[269] && f[163] && f[349] && !f[622]; // c6t126i12
	assign leaf[202] = f[269] && f[163] && f[349] && f[622]; // c6t126i12
	assign leaf[203] = !f[654] && !f[572] && !f[544] && !f[599]; // c6t136i13
	assign leaf[204] = !f[654] && !f[572] && !f[544] && f[599]; // c6t136i13
	assign leaf[205] = !f[654] && !f[572] && f[544] && !f[543]; // c6t136i13
	assign leaf[206] = !f[654] && !f[572] && f[544] && f[543]; // c6t136i13
	assign leaf[207] = !f[654] && f[572] && !f[429] && !f[431]; // c6t136i13
	assign leaf[208] = !f[654] && f[572] && !f[429] && f[431]; // c6t136i13
	assign leaf[209] = !f[654] && f[572] && f[429] && !f[593]; // c6t136i13
	assign leaf[210] = !f[654] && f[572] && f[429] && f[593]; // c6t136i13
	assign leaf[211] = f[654] && !f[132] && !f[131] && !f[164]; // c6t136i13
	assign leaf[212] = f[654] && !f[132] && !f[131] && f[164]; // c6t136i13
	assign leaf[213] = f[654] && !f[132] && f[131] && !f[430]; // c6t136i13
	assign leaf[214] = f[654] && !f[132] && f[131] && f[430]; // c6t136i13
	assign leaf[215] = f[654] && f[132] && !f[458] && !f[525]; // c6t136i13
	assign leaf[216] = f[654] && f[132] && !f[458] && f[525]; // c6t136i13
	assign leaf[217] = f[654] && f[132] && f[458] && !f[326]; // c6t136i13
	assign leaf[218] = f[654] && f[132] && f[458] && f[326]; // c6t136i13
	assign leaf[219] = !f[242] && !f[296] && !f[216] && !f[350]; // c6t146i14
	assign leaf[220] = !f[242] && !f[296] && !f[216] && f[350]; // c6t146i14
	assign leaf[221] = !f[242] && !f[296] && f[216] && !f[632]; // c6t146i14
	assign leaf[222] = !f[242] && !f[296] && f[216] && f[632]; // c6t146i14
	assign leaf[223] = !f[242] && f[296] && !f[357] && !f[131]; // c6t146i14
	assign leaf[224] = !f[242] && f[296] && !f[357] && f[131]; // c6t146i14
	assign leaf[225] = !f[242] && f[296] && f[357] && !f[485]; // c6t146i14
	assign leaf[226] = !f[242] && f[296] && f[357] && f[485]; // c6t146i14
	assign leaf[227] = f[242] && !f[164] && !f[326] && !f[131]; // c6t146i14
	assign leaf[228] = f[242] && !f[164] && !f[326] && f[131]; // c6t146i14
	assign leaf[229] = f[242] && !f[164] && f[326] && !f[387]; // c6t146i14
	assign leaf[230] = f[242] && !f[164] && f[326] && f[387]; // c6t146i14
	assign leaf[231] = f[242] && f[164] && !f[623]; // c6t146i14
	assign leaf[232] = f[242] && f[164] && f[623] && !f[622]; // c6t146i14
	assign leaf[233] = f[242] && f[164] && f[623] && f[622]; // c6t146i14
	assign leaf[234] = !f[414] && !f[430] && !f[416] && !f[431]; // c6t156i15
	assign leaf[235] = !f[414] && !f[430] && !f[416] && f[431]; // c6t156i15
	assign leaf[236] = !f[414] && !f[430] && f[416] && !f[265]; // c6t156i15
	assign leaf[237] = !f[414] && !f[430] && f[416] && f[265]; // c6t156i15
	assign leaf[238] = !f[414] && f[430] && !f[347] && !f[210]; // c6t156i15
	assign leaf[239] = !f[414] && f[430] && !f[347] && f[210]; // c6t156i15
	assign leaf[240] = !f[414] && f[430] && f[347] && !f[299]; // c6t156i15
	assign leaf[241] = !f[414] && f[430] && f[347] && f[299]; // c6t156i15
	assign leaf[242] = f[414] && !f[657] && !f[239] && !f[187]; // c6t156i15
	assign leaf[243] = f[414] && !f[657] && !f[239] && f[187]; // c6t156i15
	assign leaf[244] = f[414] && !f[657] && f[239] && !f[347]; // c6t156i15
	assign leaf[245] = f[414] && !f[657] && f[239] && f[347]; // c6t156i15
	assign leaf[246] = f[414] && f[657] && !f[454]; // c6t156i15
	assign leaf[247] = f[414] && f[657] && f[454] && !f[434]; // c6t156i15
	assign leaf[248] = f[414] && f[657] && f[454] && f[434]; // c6t156i15
	assign leaf[249] = !f[685] && !f[574] && !f[131] && !f[268]; // c6t166i16
	assign leaf[250] = !f[685] && !f[574] && !f[131] && f[268]; // c6t166i16
	assign leaf[251] = !f[685] && !f[574] && f[131] && !f[265]; // c6t166i16
	assign leaf[252] = !f[685] && !f[574] && f[131] && f[265]; // c6t166i16
	assign leaf[253] = !f[685] && f[574] && !f[210] && !f[156]; // c6t166i16
	assign leaf[254] = !f[685] && f[574] && !f[210] && f[156]; // c6t166i16
	assign leaf[255] = !f[685] && f[574] && f[210] && !f[100]; // c6t166i16
	assign leaf[256] = !f[685] && f[574] && f[210] && f[100]; // c6t166i16
	assign leaf[257] = f[685] && !f[192]; // c6t166i16
	assign leaf[258] = f[685] && f[192]; // c6t166i16
	assign leaf[259] = !f[685] && !f[623] && !f[575] && !f[269]; // c6t176i17
	assign leaf[260] = !f[685] && !f[623] && !f[575] && f[269]; // c6t176i17
	assign leaf[261] = !f[685] && !f[623] && f[575] && !f[631]; // c6t176i17
	assign leaf[262] = !f[685] && !f[623] && f[575] && f[631]; // c6t176i17
	assign leaf[263] = !f[685] && f[623] && !f[400] && !f[343]; // c6t176i17
	assign leaf[264] = !f[685] && f[623] && !f[400] && f[343]; // c6t176i17
	assign leaf[265] = !f[685] && f[623] && f[400] && !f[273]; // c6t176i17
	assign leaf[266] = !f[685] && f[623] && f[400] && f[273]; // c6t176i17
	assign leaf[267] = f[685] && !f[598]; // c6t176i17
	assign leaf[268] = f[685] && f[598] && !f[234] && !f[158]; // c6t176i17
	assign leaf[269] = f[685] && f[598] && !f[234] && f[158]; // c6t176i17
	assign leaf[270] = f[685] && f[598] && f[234]; // c6t176i17
	assign leaf[271] = !f[544] && !f[570] && !f[134] && !f[119]; // c6t186i18
	assign leaf[272] = !f[544] && !f[570] && !f[134] && f[119]; // c6t186i18
	assign leaf[273] = !f[544] && !f[570] && f[134] && !f[241]; // c6t186i18
	assign leaf[274] = !f[544] && !f[570] && f[134] && f[241]; // c6t186i18
	assign leaf[275] = !f[544] && f[570] && !f[429] && !f[291]; // c6t186i18
	assign leaf[276] = !f[544] && f[570] && !f[429] && f[291]; // c6t186i18
	assign leaf[277] = !f[544] && f[570] && f[429] && !f[160]; // c6t186i18
	assign leaf[278] = !f[544] && f[570] && f[429] && f[160]; // c6t186i18
	assign leaf[279] = f[544] && !f[653] && !f[609] && !f[296]; // c6t186i18
	assign leaf[280] = f[544] && !f[653] && !f[609] && f[296]; // c6t186i18
	assign leaf[281] = f[544] && !f[653] && f[609] && !f[455]; // c6t186i18
	assign leaf[282] = f[544] && !f[653] && f[609] && f[455]; // c6t186i18
	assign leaf[283] = f[544] && f[653] && !f[132] && !f[496]; // c6t186i18
	assign leaf[284] = f[544] && f[653] && !f[132] && f[496]; // c6t186i18
	assign leaf[285] = f[544] && f[653] && f[132] && !f[652]; // c6t186i18
	assign leaf[286] = f[544] && f[653] && f[132] && f[652]; // c6t186i18
	assign leaf[287] = !f[522] && !f[578] && !f[132] && !f[129]; // c6t196i19
	assign leaf[288] = !f[522] && !f[578] && !f[132] && f[129]; // c6t196i19
	assign leaf[289] = !f[522] && !f[578] && f[132] && !f[403]; // c6t196i19
	assign leaf[290] = !f[522] && !f[578] && f[132] && f[403]; // c6t196i19
	assign leaf[291] = !f[522] && f[578] && !f[211] && !f[400]; // c6t196i19
	assign leaf[292] = !f[522] && f[578] && !f[211] && f[400]; // c6t196i19
	assign leaf[293] = !f[522] && f[578] && f[211] && !f[234]; // c6t196i19
	assign leaf[294] = !f[522] && f[578] && f[211] && f[234]; // c6t196i19
	assign leaf[295] = f[522] && !f[207] && !f[125] && !f[622]; // c6t196i19
	assign leaf[296] = f[522] && !f[207] && !f[125] && f[622]; // c6t196i19
	assign leaf[297] = f[522] && !f[207] && f[125] && !f[236]; // c6t196i19
	assign leaf[298] = f[522] && !f[207] && f[125] && f[236]; // c6t196i19
	assign leaf[299] = f[522] && f[207] && !f[96] && !f[414]; // c6t196i19
	assign leaf[300] = f[522] && f[207] && !f[96] && f[414]; // c6t196i19
	assign leaf[301] = f[522] && f[207] && f[96] && !f[183]; // c6t196i19
	assign leaf[302] = f[522] && f[207] && f[96] && f[183]; // c6t196i19
	assign leaf[303] = !f[486] && !f[387] && !f[488] && !f[456]; // c6t206i20
	assign leaf[304] = !f[486] && !f[387] && !f[488] && f[456]; // c6t206i20
	assign leaf[305] = !f[486] && !f[387] && f[488] && !f[522]; // c6t206i20
	assign leaf[306] = !f[486] && !f[387] && f[488] && f[522]; // c6t206i20
	assign leaf[307] = !f[486] && f[387] && !f[236] && !f[291]; // c6t206i20
	assign leaf[308] = !f[486] && f[387] && !f[236] && f[291]; // c6t206i20
	assign leaf[309] = !f[486] && f[387] && f[236] && !f[356]; // c6t206i20
	assign leaf[310] = !f[486] && f[387] && f[236] && f[356]; // c6t206i20
	assign leaf[311] = f[486] && !f[430] && !f[428] && !f[485]; // c6t206i20
	assign leaf[312] = f[486] && !f[430] && !f[428] && f[485]; // c6t206i20
	assign leaf[313] = f[486] && !f[430] && f[428] && !f[212]; // c6t206i20
	assign leaf[314] = f[486] && !f[430] && f[428] && f[212]; // c6t206i20
	assign leaf[315] = f[486] && f[430] && !f[601] && !f[546]; // c6t206i20
	assign leaf[316] = f[486] && f[430] && !f[601] && f[546]; // c6t206i20
	assign leaf[317] = f[486] && f[430] && f[601] && !f[326]; // c6t206i20
	assign leaf[318] = f[486] && f[430] && f[601] && f[326]; // c6t206i20
	assign leaf[319] = !f[297] && !f[273] && !f[351] && !f[271]; // c6t216i21
	assign leaf[320] = !f[297] && !f[273] && !f[351] && f[271]; // c6t216i21
	assign leaf[321] = !f[297] && !f[273] && f[351] && !f[430]; // c6t216i21
	assign leaf[322] = !f[297] && !f[273] && f[351] && f[430]; // c6t216i21
	assign leaf[323] = !f[297] && f[273] && !f[121] && !f[328]; // c6t216i21
	assign leaf[324] = !f[297] && f[273] && !f[121] && f[328]; // c6t216i21
	assign leaf[325] = !f[297] && f[273] && f[121] && !f[326]; // c6t216i21
	assign leaf[326] = !f[297] && f[273] && f[121] && f[326]; // c6t216i21
	assign leaf[327] = f[297] && !f[329] && !f[331] && !f[384]; // c6t216i21
	assign leaf[328] = f[297] && !f[329] && !f[331] && f[384]; // c6t216i21
	assign leaf[329] = f[297] && !f[329] && f[331] && !f[245]; // c6t216i21
	assign leaf[330] = f[297] && !f[329] && f[331] && f[245]; // c6t216i21
	assign leaf[331] = f[297] && f[329] && !f[150] && !f[379]; // c6t216i21
	assign leaf[332] = f[297] && f[329] && !f[150] && f[379]; // c6t216i21
	assign leaf[333] = f[297] && f[329] && f[150] && !f[209]; // c6t216i21
	assign leaf[334] = f[297] && f[329] && f[150] && f[209]; // c6t216i21
	assign leaf[335] = !f[683] && !f[635] && !f[622] && !f[687]; // c6t226i22
	assign leaf[336] = !f[683] && !f[635] && !f[622] && f[687]; // c6t226i22
	assign leaf[337] = !f[683] && !f[635] && f[622] && !f[498]; // c6t226i22
	assign leaf[338] = !f[683] && !f[635] && f[622] && f[498]; // c6t226i22
	assign leaf[339] = !f[683] && f[635] && !f[345] && !f[518]; // c6t226i22
	assign leaf[340] = !f[683] && f[635] && !f[345] && f[518]; // c6t226i22
	assign leaf[341] = !f[683] && f[635] && f[345] && !f[245]; // c6t226i22
	assign leaf[342] = !f[683] && f[635] && f[345] && f[245]; // c6t226i22
	assign leaf[343] = f[683]; // c6t226i22
	assign leaf[344] = !f[325] && !f[301] && !f[351] && !f[299]; // c6t236i23
	assign leaf[345] = !f[325] && !f[301] && !f[351] && f[299]; // c6t236i23
	assign leaf[346] = !f[325] && !f[301] && f[351] && !f[431]; // c6t236i23
	assign leaf[347] = !f[325] && !f[301] && f[351] && f[431]; // c6t236i23
	assign leaf[348] = !f[325] && f[301] && !f[415] && !f[122]; // c6t236i23
	assign leaf[349] = !f[325] && f[301] && !f[415] && f[122]; // c6t236i23
	assign leaf[350] = !f[325] && f[301] && f[415] && !f[381]; // c6t236i23
	assign leaf[351] = !f[325] && f[301] && f[415] && f[381]; // c6t236i23
	assign leaf[352] = f[325] && !f[357] && !f[359] && !f[384]; // c6t236i23
	assign leaf[353] = f[325] && !f[357] && !f[359] && f[384]; // c6t236i23
	assign leaf[354] = f[325] && !f[357] && f[359] && !f[303]; // c6t236i23
	assign leaf[355] = f[325] && !f[357] && f[359] && f[303]; // c6t236i23
	assign leaf[356] = f[325] && f[357] && !f[268] && !f[214]; // c6t236i23
	assign leaf[357] = f[325] && f[357] && !f[268] && f[214]; // c6t236i23
	assign leaf[358] = f[325] && f[357] && f[268] && !f[490]; // c6t236i23
	assign leaf[359] = f[325] && f[357] && f[268] && f[490]; // c6t236i23
	assign leaf[360] = !f[430] && !f[399] && !f[431] && !f[387]; // c6t246i24
	assign leaf[361] = !f[430] && !f[399] && !f[431] && f[387]; // c6t246i24
	assign leaf[362] = !f[430] && !f[399] && f[431] && !f[326]; // c6t246i24
	assign leaf[363] = !f[430] && !f[399] && f[431] && f[326]; // c6t246i24
	assign leaf[364] = !f[430] && f[399] && !f[434] && !f[432]; // c6t246i24
	assign leaf[365] = !f[430] && f[399] && !f[434] && f[432]; // c6t246i24
	assign leaf[366] = !f[430] && f[399] && f[434] && !f[546]; // c6t246i24
	assign leaf[367] = !f[430] && f[399] && f[434] && f[546]; // c6t246i24
	assign leaf[368] = f[430] && !f[486] && !f[432] && !f[300]; // c6t246i24
	assign leaf[369] = f[430] && !f[486] && !f[432] && f[300]; // c6t246i24
	assign leaf[370] = f[430] && !f[486] && f[432] && !f[487]; // c6t246i24
	assign leaf[371] = f[430] && !f[486] && f[432] && f[487]; // c6t246i24
	assign leaf[372] = f[430] && f[486] && !f[374] && !f[181]; // c6t246i24
	assign leaf[373] = f[430] && f[486] && !f[374] && f[181]; // c6t246i24
	assign leaf[374] = f[430] && f[486] && f[374] && !f[571]; // c6t246i24
	assign leaf[375] = f[430] && f[486] && f[374] && f[571]; // c6t246i24
	assign leaf[376] = !f[685] && !f[325] && !f[274] && !f[351]; // c6t256i25
	assign leaf[377] = !f[685] && !f[325] && !f[274] && f[351]; // c6t256i25
	assign leaf[378] = !f[685] && !f[325] && f[274] && !f[580]; // c6t256i25
	assign leaf[379] = !f[685] && !f[325] && f[274] && f[580]; // c6t256i25
	assign leaf[380] = !f[685] && f[325] && !f[357] && !f[359]; // c6t256i25
	assign leaf[381] = !f[685] && f[325] && !f[357] && f[359]; // c6t256i25
	assign leaf[382] = !f[685] && f[325] && f[357] && !f[410]; // c6t256i25
	assign leaf[383] = !f[685] && f[325] && f[357] && f[410]; // c6t256i25
	assign leaf[384] = f[685] && !f[599]; // c6t256i25
	assign leaf[385] = f[685] && f[599] && !f[206] && !f[325]; // c6t256i25
	assign leaf[386] = f[685] && f[599] && !f[206] && f[325]; // c6t256i25
	assign leaf[387] = f[685] && f[599] && f[206]; // c6t256i25
	assign leaf[388] = !f[683] && !f[609] && !f[403] && !f[414]; // c6t266i26
	assign leaf[389] = !f[683] && !f[609] && !f[403] && f[414]; // c6t266i26
	assign leaf[390] = !f[683] && !f[609] && f[403] && !f[487]; // c6t266i26
	assign leaf[391] = !f[683] && !f[609] && f[403] && f[487]; // c6t266i26
	assign leaf[392] = !f[683] && f[609] && !f[455] && !f[487]; // c6t266i26
	assign leaf[393] = !f[683] && f[609] && !f[455] && f[487]; // c6t266i26
	assign leaf[394] = !f[683] && f[609] && f[455] && !f[638]; // c6t266i26
	assign leaf[395] = !f[683] && f[609] && f[455] && f[638]; // c6t266i26
	assign leaf[396] = f[683]; // c6t266i26
	assign leaf[397] = !f[209] && !f[154] && !f[575] && !f[520]; // c6t276i27
	assign leaf[398] = !f[209] && !f[154] && !f[575] && f[520]; // c6t276i27
	assign leaf[399] = !f[209] && !f[154] && f[575] && !f[291]; // c6t276i27
	assign leaf[400] = !f[209] && !f[154] && f[575] && f[291]; // c6t276i27
	assign leaf[401] = !f[209] && f[154] && !f[416] && !f[183]; // c6t276i27
	assign leaf[402] = !f[209] && f[154] && !f[416] && f[183]; // c6t276i27
	assign leaf[403] = !f[209] && f[154] && f[416] && !f[383]; // c6t276i27
	assign leaf[404] = !f[209] && f[154] && f[416] && f[383]; // c6t276i27
	assign leaf[405] = f[209] && !f[128] && !f[99] && !f[130]; // c6t276i27
	assign leaf[406] = f[209] && !f[128] && !f[99] && f[130]; // c6t276i27
	assign leaf[407] = f[209] && !f[128] && f[99] && !f[410]; // c6t276i27
	assign leaf[408] = f[209] && !f[128] && f[99] && f[410]; // c6t276i27
	assign leaf[409] = f[209] && f[128] && !f[430] && !f[351]; // c6t276i27
	assign leaf[410] = f[209] && f[128] && !f[430] && f[351]; // c6t276i27
	assign leaf[411] = f[209] && f[128] && f[430] && !f[292]; // c6t276i27
	assign leaf[412] = f[209] && f[128] && f[430] && f[292]; // c6t276i27
	assign leaf[413] = !f[686] && !f[623] && !f[163] && !f[269]; // c6t286i28
	assign leaf[414] = !f[686] && !f[623] && !f[163] && f[269]; // c6t286i28
	assign leaf[415] = !f[686] && !f[623] && f[163] && !f[597]; // c6t286i28
	assign leaf[416] = !f[686] && !f[623] && f[163] && f[597]; // c6t286i28
	assign leaf[417] = !f[686] && f[623] && !f[400] && !f[599]; // c6t286i28
	assign leaf[418] = !f[686] && f[623] && !f[400] && f[599]; // c6t286i28
	assign leaf[419] = !f[686] && f[623] && f[400] && !f[511]; // c6t286i28
	assign leaf[420] = !f[686] && f[623] && f[400] && f[511]; // c6t286i28
	assign leaf[421] = f[686] && !f[569]; // c6t286i28
	assign leaf[422] = f[686] && f[569] && !f[234]; // c6t286i28
	assign leaf[423] = f[686] && f[569] && f[234]; // c6t286i28
	assign leaf[424] = !f[652] && !f[544] && !f[570] && !f[569]; // c6t296i29
	assign leaf[425] = !f[652] && !f[544] && !f[570] && f[569]; // c6t296i29
	assign leaf[426] = !f[652] && !f[544] && f[570] && !f[428]; // c6t296i29
	assign leaf[427] = !f[652] && !f[544] && f[570] && f[428]; // c6t296i29
	assign leaf[428] = !f[652] && f[544] && !f[236] && !f[153]; // c6t296i29
	assign leaf[429] = !f[652] && f[544] && !f[236] && f[153]; // c6t296i29
	assign leaf[430] = !f[652] && f[544] && f[236] && !f[322]; // c6t296i29
	assign leaf[431] = !f[652] && f[544] && f[236] && f[322]; // c6t296i29
	assign leaf[432] = f[652] && !f[133] && !f[498]; // c6t296i29
	assign leaf[433] = f[652] && !f[133] && f[498]; // c6t296i29
	assign leaf[434] = f[652] && f[133] && !f[292]; // c6t296i29
	assign leaf[435] = f[652] && f[133] && f[292]; // c6t296i29
	assign leaf[436] = !f[684] && !f[622] && !f[163] && !f[516]; // c6t306i30
	assign leaf[437] = !f[684] && !f[622] && !f[163] && f[516]; // c6t306i30
	assign leaf[438] = !f[684] && !f[622] && f[163] && !f[324]; // c6t306i30
	assign leaf[439] = !f[684] && !f[622] && f[163] && f[324]; // c6t306i30
	assign leaf[440] = !f[684] && f[622] && !f[498]; // c6t306i30
	assign leaf[441] = !f[684] && f[622] && f[498]; // c6t306i30
	assign leaf[442] = f[684] && !f[408] && !f[572]; // c6t306i30
	assign leaf[443] = f[684] && !f[408] && f[572]; // c6t306i30
	assign leaf[444] = f[684] && f[408]; // c6t306i30
	assign leaf[445] = !f[602] && !f[547] && !f[630] && !f[164]; // c6t316i31
	assign leaf[446] = !f[602] && !f[547] && !f[630] && f[164]; // c6t316i31
	assign leaf[447] = !f[602] && !f[547] && f[630] && !f[206]; // c6t316i31
	assign leaf[448] = !f[602] && !f[547] && f[630] && f[206]; // c6t316i31
	assign leaf[449] = !f[602] && f[547] && !f[236] && !f[155]; // c6t316i31
	assign leaf[450] = !f[602] && f[547] && !f[236] && f[155]; // c6t316i31
	assign leaf[451] = !f[602] && f[547] && f[236] && !f[383]; // c6t316i31
	assign leaf[452] = !f[602] && f[547] && f[236] && f[383]; // c6t316i31
	assign leaf[453] = f[602] && !f[400] && !f[459] && !f[359]; // c6t316i31
	assign leaf[454] = f[602] && !f[400] && !f[459] && f[359]; // c6t316i31
	assign leaf[455] = f[602] && !f[400] && f[459] && !f[326]; // c6t316i31
	assign leaf[456] = f[602] && !f[400] && f[459] && f[326]; // c6t316i31
	assign leaf[457] = f[602] && f[400] && !f[382] && !f[483]; // c6t316i31
	assign leaf[458] = f[602] && f[400] && !f[382] && f[483]; // c6t316i31
	assign leaf[459] = f[602] && f[400] && f[382] && !f[441]; // c6t316i31
	assign leaf[460] = f[602] && f[400] && f[382] && f[441]; // c6t316i31
	assign leaf[461] = !f[522] && !f[409] && !f[519] && !f[525]; // c6t326i32
	assign leaf[462] = !f[522] && !f[409] && !f[519] && f[525]; // c6t326i32
	assign leaf[463] = !f[522] && !f[409] && f[519] && !f[209]; // c6t326i32
	assign leaf[464] = !f[522] && !f[409] && f[519] && f[209]; // c6t326i32
	assign leaf[465] = !f[522] && f[409] && !f[525] && !f[319]; // c6t326i32
	assign leaf[466] = !f[522] && f[409] && !f[525] && f[319]; // c6t326i32
	assign leaf[467] = !f[522] && f[409] && f[525] && !f[322]; // c6t326i32
	assign leaf[468] = !f[522] && f[409] && f[525] && f[322]; // c6t326i32
	assign leaf[469] = f[522] && !f[402] && !f[387] && !f[212]; // c6t326i32
	assign leaf[470] = f[522] && !f[402] && !f[387] && f[212]; // c6t326i32
	assign leaf[471] = f[522] && !f[402] && f[387] && !f[264]; // c6t326i32
	assign leaf[472] = f[522] && !f[402] && f[387] && f[264]; // c6t326i32
	assign leaf[473] = f[522] && f[402] && !f[178] && !f[301]; // c6t326i32
	assign leaf[474] = f[522] && f[402] && !f[178] && f[301]; // c6t326i32
	assign leaf[475] = f[522] && f[402] && f[178] && !f[210]; // c6t326i32
	assign leaf[476] = f[522] && f[402] && f[178] && f[210]; // c6t326i32
	assign leaf[477] = !f[683] && !f[459] && !f[457] && !f[454]; // c6t336i33
	assign leaf[478] = !f[683] && !f[459] && !f[457] && f[454]; // c6t336i33
	assign leaf[479] = !f[683] && !f[459] && f[457] && !f[462]; // c6t336i33
	assign leaf[480] = !f[683] && !f[459] && f[457] && f[462]; // c6t336i33
	assign leaf[481] = !f[683] && f[459] && !f[375] && !f[292]; // c6t336i33
	assign leaf[482] = !f[683] && f[459] && !f[375] && f[292]; // c6t336i33
	assign leaf[483] = !f[683] && f[459] && f[375] && !f[303]; // c6t336i33
	assign leaf[484] = !f[683] && f[459] && f[375] && f[303]; // c6t336i33
	assign leaf[485] = f[683]; // c6t336i33
	assign leaf[486] = !f[683] && !f[234] && !f[151] && !f[326]; // c6t346i34
	assign leaf[487] = !f[683] && !f[234] && !f[151] && f[326]; // c6t346i34
	assign leaf[488] = !f[683] && !f[234] && f[151] && !f[398]; // c6t346i34
	assign leaf[489] = !f[683] && !f[234] && f[151] && f[398]; // c6t346i34
	assign leaf[490] = !f[683] && f[234] && !f[266] && !f[545]; // c6t346i34
	assign leaf[491] = !f[683] && f[234] && !f[266] && f[545]; // c6t346i34
	assign leaf[492] = !f[683] && f[234] && f[266] && !f[272]; // c6t346i34
	assign leaf[493] = !f[683] && f[234] && f[266] && f[272]; // c6t346i34
	assign leaf[494] = f[683]; // c6t346i34
	assign leaf[495] = !f[601] && !f[64] && !f[295] && !f[241]; // c6t356i35
	assign leaf[496] = !f[601] && !f[64] && !f[295] && f[241]; // c6t356i35
	assign leaf[497] = !f[601] && !f[64] && f[295] && !f[132]; // c6t356i35
	assign leaf[498] = !f[601] && !f[64] && f[295] && f[132]; // c6t356i35
	assign leaf[499] = !f[601] && f[64]; // c6t356i35
	assign leaf[500] = f[601] && !f[486] && !f[455] && !f[516]; // c6t356i35
	assign leaf[501] = f[601] && !f[486] && !f[455] && f[516]; // c6t356i35
	assign leaf[502] = f[601] && !f[486] && f[455] && !f[370]; // c6t356i35
	assign leaf[503] = f[601] && !f[486] && f[455] && f[370]; // c6t356i35
	assign leaf[504] = f[601] && f[486] && !f[374] && !f[181]; // c6t356i35
	assign leaf[505] = f[601] && f[486] && !f[374] && f[181]; // c6t356i35
	assign leaf[506] = f[601] && f[486] && f[374] && !f[458]; // c6t356i35
	assign leaf[507] = f[601] && f[486] && f[374] && f[458]; // c6t356i35
	assign leaf[508] = !f[637] && !f[299] && !f[301] && !f[324]; // c6t366i36
	assign leaf[509] = !f[637] && !f[299] && !f[301] && f[324]; // c6t366i36
	assign leaf[510] = !f[637] && !f[299] && f[301] && !f[122]; // c6t366i36
	assign leaf[511] = !f[637] && !f[299] && f[301] && f[122]; // c6t366i36
	assign leaf[512] = !f[637] && f[299] && !f[382] && !f[176]; // c6t366i36
	assign leaf[513] = !f[637] && f[299] && !f[382] && f[176]; // c6t366i36
	assign leaf[514] = !f[637] && f[299] && f[382] && !f[357]; // c6t366i36
	assign leaf[515] = !f[637] && f[299] && f[382] && f[357]; // c6t366i36
	assign leaf[516] = f[637] && !f[511] && !f[526] && !f[125]; // c6t366i36
	assign leaf[517] = f[637] && !f[511] && !f[526] && f[125]; // c6t366i36
	assign leaf[518] = f[637] && !f[511] && f[526]; // c6t366i36
	assign leaf[519] = f[637] && f[511] && !f[263]; // c6t366i36
	assign leaf[520] = f[637] && f[511] && f[263]; // c6t366i36
	assign leaf[521] = !f[653] && !f[689] && !f[517] && !f[151]; // c6t376i37
	assign leaf[522] = !f[653] && !f[689] && !f[517] && f[151]; // c6t376i37
	assign leaf[523] = !f[653] && !f[689] && f[517] && !f[240]; // c6t376i37
	assign leaf[524] = !f[653] && !f[689] && f[517] && f[240]; // c6t376i37
	assign leaf[525] = !f[653] && f[689] && !f[598]; // c6t376i37
	assign leaf[526] = !f[653] && f[689] && f[598]; // c6t376i37
	assign leaf[527] = f[653] && !f[162] && !f[627] && !f[519]; // c6t376i37
	assign leaf[528] = f[653] && !f[162] && !f[627] && f[519]; // c6t376i37
	assign leaf[529] = f[653] && !f[162] && f[627]; // c6t376i37
	assign leaf[530] = f[653] && f[162] && !f[490] && !f[539]; // c6t376i37
	assign leaf[531] = f[653] && f[162] && !f[490] && f[539]; // c6t376i37
	assign leaf[532] = f[653] && f[162] && f[490]; // c6t376i37
	assign leaf[533] = !f[622] && !f[159] && !f[239] && !f[574]; // c6t386i38
	assign leaf[534] = !f[622] && !f[159] && !f[239] && f[574]; // c6t386i38
	assign leaf[535] = !f[622] && !f[159] && f[239] && !f[156]; // c6t386i38
	assign leaf[536] = !f[622] && !f[159] && f[239] && f[156]; // c6t386i38
	assign leaf[537] = !f[622] && f[159] && !f[325] && !f[328]; // c6t386i38
	assign leaf[538] = !f[622] && f[159] && !f[325] && f[328]; // c6t386i38
	assign leaf[539] = !f[622] && f[159] && f[325] && !f[467]; // c6t386i38
	assign leaf[540] = !f[622] && f[159] && f[325] && f[467]; // c6t386i38
	assign leaf[541] = f[622]; // c6t386i38
	assign leaf[542] = !f[91] && !f[682] && !f[459] && !f[457]; // c6t396i39
	assign leaf[543] = !f[91] && !f[682] && !f[459] && f[457]; // c6t396i39
	assign leaf[544] = !f[91] && !f[682] && f[459] && !f[403]; // c6t396i39
	assign leaf[545] = !f[91] && !f[682] && f[459] && f[403]; // c6t396i39
	assign leaf[546] = !f[91] && f[682]; // c6t396i39
	assign leaf[547] = f[91] && !f[356]; // c6t396i39
	assign leaf[548] = f[91] && f[356]; // c6t396i39
	assign leaf[549] = !f[609] && !f[93] && !f[270] && !f[274]; // c6t406i40
	assign leaf[550] = !f[609] && !f[93] && !f[270] && f[274]; // c6t406i40
	assign leaf[551] = !f[609] && !f[93] && f[270] && !f[350]; // c6t406i40
	assign leaf[552] = !f[609] && !f[93] && f[270] && f[350]; // c6t406i40
	assign leaf[553] = !f[609] && f[93] && !f[123] && !f[431]; // c6t406i40
	assign leaf[554] = !f[609] && f[93] && !f[123] && f[431]; // c6t406i40
	assign leaf[555] = !f[609] && f[93] && f[123] && !f[206]; // c6t406i40
	assign leaf[556] = !f[609] && f[93] && f[123] && f[206]; // c6t406i40
	assign leaf[557] = f[609] && !f[455] && !f[551] && !f[290]; // c6t406i40
	assign leaf[558] = f[609] && !f[455] && !f[551] && f[290]; // c6t406i40
	assign leaf[559] = f[609] && !f[455] && f[551] && !f[555]; // c6t406i40
	assign leaf[560] = f[609] && !f[455] && f[551] && f[555]; // c6t406i40
	assign leaf[561] = f[609] && f[455] && !f[633] && !f[573]; // c6t406i40
	assign leaf[562] = f[609] && f[455] && !f[633] && f[573]; // c6t406i40
	assign leaf[563] = f[609] && f[455] && f[633] && !f[205]; // c6t406i40
	assign leaf[564] = f[609] && f[455] && f[633] && f[205]; // c6t406i40
	assign leaf[565] = !f[622] && !f[208] && !f[98] && !f[550]; // c6t416i41
	assign leaf[566] = !f[622] && !f[208] && !f[98] && f[550]; // c6t416i41
	assign leaf[567] = !f[622] && !f[208] && f[98] && !f[551]; // c6t416i41
	assign leaf[568] = !f[622] && !f[208] && f[98] && f[551]; // c6t416i41
	assign leaf[569] = !f[622] && f[208] && !f[318] && !f[416]; // c6t416i41
	assign leaf[570] = !f[622] && f[208] && !f[318] && f[416]; // c6t416i41
	assign leaf[571] = !f[622] && f[208] && f[318] && !f[178]; // c6t416i41
	assign leaf[572] = !f[622] && f[208] && f[318] && f[178]; // c6t416i41
	assign leaf[573] = f[622]; // c6t416i41
	assign leaf[574] = !f[594] && !f[685] && !f[661] && !f[635]; // c6t426i42
	assign leaf[575] = !f[594] && !f[685] && !f[661] && f[635]; // c6t426i42
	assign leaf[576] = !f[594] && !f[685] && f[661] && !f[158]; // c6t426i42
	assign leaf[577] = !f[594] && !f[685] && f[661] && f[158]; // c6t426i42
	assign leaf[578] = !f[594] && f[685] && !f[598]; // c6t426i42
	assign leaf[579] = !f[594] && f[685] && f[598] && !f[381]; // c6t426i42
	assign leaf[580] = !f[594] && f[685] && f[598] && f[381]; // c6t426i42
	assign leaf[581] = f[594] && !f[400] && !f[185] && !f[543]; // c6t426i42
	assign leaf[582] = f[594] && !f[400] && !f[185] && f[543]; // c6t426i42
	assign leaf[583] = f[594] && !f[400] && f[185]; // c6t426i42
	assign leaf[584] = f[594] && f[400] && !f[217] && !f[435]; // c6t426i42
	assign leaf[585] = f[594] && f[400] && !f[217] && f[435]; // c6t426i42
	assign leaf[586] = f[594] && f[400] && f[217]; // c6t426i42
	assign leaf[587] = !f[275] && !f[101] && !f[163] && !f[268]; // c6t436i43
	assign leaf[588] = !f[275] && !f[101] && !f[163] && f[268]; // c6t436i43
	assign leaf[589] = !f[275] && !f[101] && f[163] && !f[355]; // c6t436i43
	assign leaf[590] = !f[275] && !f[101] && f[163] && f[355]; // c6t436i43
	assign leaf[591] = !f[275] && f[101] && !f[74] && !f[547]; // c6t436i43
	assign leaf[592] = !f[275] && f[101] && !f[74] && f[547]; // c6t436i43
	assign leaf[593] = !f[275] && f[101] && f[74] && !f[485]; // c6t436i43
	assign leaf[594] = !f[275] && f[101] && f[74] && f[485]; // c6t436i43
	assign leaf[595] = f[275] && !f[272]; // c6t436i43
	assign leaf[596] = f[275] && f[272] && !f[332] && !f[515]; // c6t436i43
	assign leaf[597] = f[275] && f[272] && !f[332] && f[515]; // c6t436i43
	assign leaf[598] = f[275] && f[272] && f[332]; // c6t436i43
	assign leaf[599] = !f[517] && !f[178] && !f[600] && !f[317]; // c6t446i44
	assign leaf[600] = !f[517] && !f[178] && !f[600] && f[317]; // c6t446i44
	assign leaf[601] = !f[517] && !f[178] && f[600] && !f[574]; // c6t446i44
	assign leaf[602] = !f[517] && !f[178] && f[600] && f[574]; // c6t446i44
	assign leaf[603] = !f[517] && f[178] && !f[319] && !f[184]; // c6t446i44
	assign leaf[604] = !f[517] && f[178] && !f[319] && f[184]; // c6t446i44
	assign leaf[605] = !f[517] && f[178] && f[319] && !f[428]; // c6t446i44
	assign leaf[606] = !f[517] && f[178] && f[319] && f[428]; // c6t446i44
	assign leaf[607] = f[517] && !f[652] && !f[602] && !f[383]; // c6t446i44
	assign leaf[608] = f[517] && !f[652] && !f[602] && f[383]; // c6t446i44
	assign leaf[609] = f[517] && !f[652] && f[602] && !f[381]; // c6t446i44
	assign leaf[610] = f[517] && !f[652] && f[602] && f[381]; // c6t446i44
	assign leaf[611] = f[517] && f[652]; // c6t446i44
	assign leaf[612] = !f[682] && !f[459] && !f[387] && !f[429]; // c6t456i45
	assign leaf[613] = !f[682] && !f[459] && !f[387] && f[429]; // c6t456i45
	assign leaf[614] = !f[682] && !f[459] && f[387] && !f[409]; // c6t456i45
	assign leaf[615] = !f[682] && !f[459] && f[387] && f[409]; // c6t456i45
	assign leaf[616] = !f[682] && f[459] && !f[544] && !f[159]; // c6t456i45
	assign leaf[617] = !f[682] && f[459] && !f[544] && f[159]; // c6t456i45
	assign leaf[618] = !f[682] && f[459] && f[544] && !f[487]; // c6t456i45
	assign leaf[619] = !f[682] && f[459] && f[544] && f[487]; // c6t456i45
	assign leaf[620] = f[682]; // c6t456i45
	assign leaf[621] = !f[622] && !f[132] && !f[267] && !f[213]; // c6t466i46
	assign leaf[622] = !f[622] && !f[132] && !f[267] && f[213]; // c6t466i46
	assign leaf[623] = !f[622] && !f[132] && f[267] && !f[263]; // c6t466i46
	assign leaf[624] = !f[622] && !f[132] && f[267] && f[263]; // c6t466i46
	assign leaf[625] = !f[622] && f[132] && !f[326] && !f[233]; // c6t466i46
	assign leaf[626] = !f[622] && f[132] && !f[326] && f[233]; // c6t466i46
	assign leaf[627] = !f[622] && f[132] && f[326] && !f[496]; // c6t466i46
	assign leaf[628] = !f[622] && f[132] && f[326] && f[496]; // c6t466i46
	assign leaf[629] = f[622]; // c6t466i46
	assign leaf[630] = !f[455] && !f[596] && !f[607] && !f[661]; // c6t476i47
	assign leaf[631] = !f[455] && !f[596] && !f[607] && f[661]; // c6t476i47
	assign leaf[632] = !f[455] && !f[596] && f[607] && !f[457]; // c6t476i47
	assign leaf[633] = !f[455] && !f[596] && f[607] && f[457]; // c6t476i47
	assign leaf[634] = !f[455] && f[596] && !f[370] && !f[457]; // c6t476i47
	assign leaf[635] = !f[455] && f[596] && !f[370] && f[457]; // c6t476i47
	assign leaf[636] = !f[455] && f[596] && f[370]; // c6t476i47
	assign leaf[637] = f[455] && !f[601] && !f[275] && !f[546]; // c6t476i47
	assign leaf[638] = f[455] && !f[601] && !f[275] && f[546]; // c6t476i47
	assign leaf[639] = f[455] && !f[601] && f[275]; // c6t476i47
	assign leaf[640] = f[455] && f[601] && !f[186] && !f[238]; // c6t476i47
	assign leaf[641] = f[455] && f[601] && !f[186] && f[238]; // c6t476i47
	assign leaf[642] = f[455] && f[601] && f[186] && !f[346]; // c6t476i47
	assign leaf[643] = f[455] && f[601] && f[186] && f[346]; // c6t476i47
	assign leaf[644] = !f[163] && !f[269] && !f[295] && !f[185]; // c6t486i48
	assign leaf[645] = !f[163] && !f[269] && !f[295] && f[185]; // c6t486i48
	assign leaf[646] = !f[163] && !f[269] && f[295] && !f[185]; // c6t486i48
	assign leaf[647] = !f[163] && !f[269] && f[295] && f[185]; // c6t486i48
	assign leaf[648] = !f[163] && f[269] && !f[350] && !f[525]; // c6t486i48
	assign leaf[649] = !f[163] && f[269] && !f[350] && f[525]; // c6t486i48
	assign leaf[650] = !f[163] && f[269] && f[350] && !f[380]; // c6t486i48
	assign leaf[651] = !f[163] && f[269] && f[350] && f[380]; // c6t486i48
	assign leaf[652] = f[163] && !f[328] && !f[492] && !f[515]; // c6t486i48
	assign leaf[653] = f[163] && !f[328] && !f[492] && f[515]; // c6t486i48
	assign leaf[654] = f[163] && !f[328] && f[492] && !f[220]; // c6t486i48
	assign leaf[655] = f[163] && !f[328] && f[492] && f[220]; // c6t486i48
	assign leaf[656] = f[163] && f[328]; // c6t486i48
	assign leaf[657] = !f[299] && !f[301] && !f[245] && !f[324]; // c6t496i49
	assign leaf[658] = !f[299] && !f[301] && !f[245] && f[324]; // c6t496i49
	assign leaf[659] = !f[299] && !f[301] && f[245] && !f[541]; // c6t496i49
	assign leaf[660] = !f[299] && !f[301] && f[245] && f[541]; // c6t496i49
	assign leaf[661] = !f[299] && f[301] && !f[260]; // c6t496i49
	assign leaf[662] = !f[299] && f[301] && f[260] && !f[358]; // c6t496i49
	assign leaf[663] = !f[299] && f[301] && f[260] && f[358]; // c6t496i49
	assign leaf[664] = f[299] && !f[382] && !f[512] && !f[149]; // c6t496i49
	assign leaf[665] = f[299] && !f[382] && !f[512] && f[149]; // c6t496i49
	assign leaf[666] = f[299] && !f[382] && f[512] && !f[571]; // c6t496i49
	assign leaf[667] = f[299] && !f[382] && f[512] && f[571]; // c6t496i49
	assign leaf[668] = f[299] && f[382] && !f[357] && !f[456]; // c6t496i49
	assign leaf[669] = f[299] && f[382] && !f[357] && f[456]; // c6t496i49
	assign leaf[670] = f[299] && f[382] && f[357] && !f[383]; // c6t496i49
	assign leaf[671] = f[299] && f[382] && f[357] && f[383]; // c6t496i49
	assign leaf[672] = !f[652] && !f[160] && !f[240] && !f[213]; // c6t506i50
	assign leaf[673] = !f[652] && !f[160] && !f[240] && f[213]; // c6t506i50
	assign leaf[674] = !f[652] && !f[160] && f[240] && !f[158]; // c6t506i50
	assign leaf[675] = !f[652] && !f[160] && f[240] && f[158]; // c6t506i50
	assign leaf[676] = !f[652] && f[160] && !f[274] && !f[353]; // c6t506i50
	assign leaf[677] = !f[652] && f[160] && !f[274] && f[353]; // c6t506i50
	assign leaf[678] = !f[652] && f[160] && f[274]; // c6t506i50
	assign leaf[679] = f[652] && !f[163]; // c6t506i50
	assign leaf[680] = f[652] && f[163]; // c6t506i50
	assign leaf[681] = !f[428] && !f[235] && !f[124] && !f[567]; // c6t516i51
	assign leaf[682] = !f[428] && !f[235] && !f[124] && f[567]; // c6t516i51
	assign leaf[683] = !f[428] && !f[235] && f[124] && !f[426]; // c6t516i51
	assign leaf[684] = !f[428] && !f[235] && f[124] && f[426]; // c6t516i51
	assign leaf[685] = !f[428] && f[235] && !f[96] && !f[98]; // c6t516i51
	assign leaf[686] = !f[428] && f[235] && !f[96] && f[98]; // c6t516i51
	assign leaf[687] = !f[428] && f[235] && f[96] && !f[599]; // c6t516i51
	assign leaf[688] = !f[428] && f[235] && f[96] && f[599]; // c6t516i51
	assign leaf[689] = f[428] && !f[541] && !f[236] && !f[548]; // c6t516i51
	assign leaf[690] = f[428] && !f[541] && !f[236] && f[548]; // c6t516i51
	assign leaf[691] = f[428] && !f[541] && f[236] && !f[151]; // c6t516i51
	assign leaf[692] = f[428] && !f[541] && f[236] && f[151]; // c6t516i51
	assign leaf[693] = f[428] && f[541] && !f[318] && !f[264]; // c6t516i51
	assign leaf[694] = f[428] && f[541] && !f[318] && f[264]; // c6t516i51
	assign leaf[695] = f[428] && f[541] && f[318] && !f[157]; // c6t516i51
	assign leaf[696] = f[428] && f[541] && f[318] && f[157]; // c6t516i51
	assign leaf[697] = !f[409] && !f[98] && !f[571] && !f[323]; // c6t526i52
	assign leaf[698] = !f[409] && !f[98] && !f[571] && f[323]; // c6t526i52
	assign leaf[699] = !f[409] && !f[98] && f[571] && !f[271]; // c6t526i52
	assign leaf[700] = !f[409] && !f[98] && f[571] && f[271]; // c6t526i52
	assign leaf[701] = !f[409] && f[98] && !f[579] && !f[353]; // c6t526i52
	assign leaf[702] = !f[409] && f[98] && !f[579] && f[353]; // c6t526i52
	assign leaf[703] = !f[409] && f[98] && f[579] && !f[601]; // c6t526i52
	assign leaf[704] = !f[409] && f[98] && f[579] && f[601]; // c6t526i52
	assign leaf[705] = f[409] && !f[441] && !f[327] && !f[325]; // c6t526i52
	assign leaf[706] = f[409] && !f[441] && !f[327] && f[325]; // c6t526i52
	assign leaf[707] = f[409] && !f[441] && f[327] && !f[149]; // c6t526i52
	assign leaf[708] = f[409] && !f[441] && f[327] && f[149]; // c6t526i52
	assign leaf[709] = f[409] && f[441] && !f[377] && !f[270]; // c6t526i52
	assign leaf[710] = f[409] && f[441] && !f[377] && f[270]; // c6t526i52
	assign leaf[711] = f[409] && f[441] && f[377] && !f[484]; // c6t526i52
	assign leaf[712] = f[409] && f[441] && f[377] && f[484]; // c6t526i52
	assign leaf[713] = !f[91] && !f[202] && !f[439] && !f[409]; // c6t536i53
	assign leaf[714] = !f[91] && !f[202] && !f[439] && f[409]; // c6t536i53
	assign leaf[715] = !f[91] && !f[202] && f[439] && !f[403]; // c6t536i53
	assign leaf[716] = !f[91] && !f[202] && f[439] && f[403]; // c6t536i53
	assign leaf[717] = !f[91] && f[202] && !f[426]; // c6t536i53
	assign leaf[718] = !f[91] && f[202] && f[426]; // c6t536i53
	assign leaf[719] = f[91]; // c6t536i53
	assign leaf[720] = !f[295] && !f[214] && !f[635] && !f[627]; // c6t546i54
	assign leaf[721] = !f[295] && !f[214] && !f[635] && f[627]; // c6t546i54
	assign leaf[722] = !f[295] && !f[214] && f[635] && !f[130]; // c6t546i54
	assign leaf[723] = !f[295] && !f[214] && f[635] && f[130]; // c6t546i54
	assign leaf[724] = !f[295] && f[214] && !f[663] && !f[657]; // c6t546i54
	assign leaf[725] = !f[295] && f[214] && !f[663] && f[657]; // c6t546i54
	assign leaf[726] = !f[295] && f[214] && f[663]; // c6t546i54
	assign leaf[727] = f[295] && !f[237] && !f[291] && !f[321]; // c6t546i54
	assign leaf[728] = f[295] && !f[237] && !f[291] && f[321]; // c6t546i54
	assign leaf[729] = f[295] && !f[237] && f[291] && !f[207]; // c6t546i54
	assign leaf[730] = f[295] && !f[237] && f[291] && f[207]; // c6t546i54
	assign leaf[731] = f[295] && f[237] && !f[374] && !f[323]; // c6t546i54
	assign leaf[732] = f[295] && f[237] && !f[374] && f[323]; // c6t546i54
	assign leaf[733] = f[295] && f[237] && f[374] && !f[155]; // c6t546i54
	assign leaf[734] = f[295] && f[237] && f[374] && f[155]; // c6t546i54
	assign leaf[735] = !f[639] && !f[517] && !f[512] && !f[407]; // c6t556i55
	assign leaf[736] = !f[639] && !f[517] && !f[512] && f[407]; // c6t556i55
	assign leaf[737] = !f[639] && !f[517] && f[512] && !f[373]; // c6t556i55
	assign leaf[738] = !f[639] && !f[517] && f[512] && f[373]; // c6t556i55
	assign leaf[739] = !f[639] && f[517] && !f[574] && !f[515]; // c6t556i55
	assign leaf[740] = !f[639] && f[517] && !f[574] && f[515]; // c6t556i55
	assign leaf[741] = !f[639] && f[517] && f[574] && !f[239]; // c6t556i55
	assign leaf[742] = !f[639] && f[517] && f[574] && f[239]; // c6t556i55
	assign leaf[743] = f[639]; // c6t556i55
	assign leaf[744] = !f[684] && !f[302] && !f[455] && !f[288]; // c6t566i56
	assign leaf[745] = !f[684] && !f[302] && !f[455] && f[288]; // c6t566i56
	assign leaf[746] = !f[684] && !f[302] && f[455] && !f[511]; // c6t566i56
	assign leaf[747] = !f[684] && !f[302] && f[455] && f[511]; // c6t566i56
	assign leaf[748] = !f[684] && f[302] && !f[402] && !f[298]; // c6t566i56
	assign leaf[749] = !f[684] && f[302] && !f[402] && f[298]; // c6t566i56
	assign leaf[750] = !f[684] && f[302] && f[402] && !f[127]; // c6t566i56
	assign leaf[751] = !f[684] && f[302] && f[402] && f[127]; // c6t566i56
	assign leaf[752] = f[684] && !f[513]; // c6t566i56
	assign leaf[753] = f[684] && f[513]; // c6t566i56
	assign leaf[754] = !f[495] && !f[494] && !f[497] && !f[131]; // c6t576i57
	assign leaf[755] = !f[495] && !f[494] && !f[497] && f[131]; // c6t576i57
	assign leaf[756] = !f[495] && !f[494] && f[497] && !f[348]; // c6t576i57
	assign leaf[757] = !f[495] && !f[494] && f[497] && f[348]; // c6t576i57
	assign leaf[758] = !f[495] && f[494] && !f[234] && !f[544]; // c6t576i57
	assign leaf[759] = !f[495] && f[494] && !f[234] && f[544]; // c6t576i57
	assign leaf[760] = !f[495] && f[494] && f[234] && !f[439]; // c6t576i57
	assign leaf[761] = !f[495] && f[494] && f[234] && f[439]; // c6t576i57
	assign leaf[762] = f[495] && !f[431] && !f[464] && !f[434]; // c6t576i57
	assign leaf[763] = f[495] && !f[431] && !f[464] && f[434]; // c6t576i57
	assign leaf[764] = f[495] && !f[431] && f[464] && !f[487]; // c6t576i57
	assign leaf[765] = f[495] && !f[431] && f[464] && f[487]; // c6t576i57
	assign leaf[766] = f[495] && f[431] && !f[230] && !f[302]; // c6t576i57
	assign leaf[767] = f[495] && f[431] && !f[230] && f[302]; // c6t576i57
	assign leaf[768] = f[495] && f[431] && f[230]; // c6t576i57
	assign leaf[769] = !f[101] && !f[72] && !f[684] && !f[602]; // c6t586i58
	assign leaf[770] = !f[101] && !f[72] && !f[684] && f[602]; // c6t586i58
	assign leaf[771] = !f[101] && !f[72] && f[684] && !f[570]; // c6t586i58
	assign leaf[772] = !f[101] && !f[72] && f[684] && f[570]; // c6t586i58
	assign leaf[773] = !f[101] && f[72]; // c6t586i58
	assign leaf[774] = f[101] && !f[293] && !f[521] && !f[209]; // c6t586i58
	assign leaf[775] = f[101] && !f[293] && !f[521] && f[209]; // c6t586i58
	assign leaf[776] = f[101] && !f[293] && f[521] && !f[463]; // c6t586i58
	assign leaf[777] = f[101] && !f[293] && f[521] && f[463]; // c6t586i58
	assign leaf[778] = f[101] && f[293] && !f[126] && !f[544]; // c6t586i58
	assign leaf[779] = f[101] && f[293] && !f[126] && f[544]; // c6t586i58
	assign leaf[780] = f[101] && f[293] && f[126] && !f[626]; // c6t586i58
	assign leaf[781] = f[101] && f[293] && f[126] && f[626]; // c6t586i58
	assign leaf[782] = !f[601] && !f[164] && !f[128] && !f[547]; // c6t596i59
	assign leaf[783] = !f[601] && !f[164] && !f[128] && f[547]; // c6t596i59
	assign leaf[784] = !f[601] && !f[164] && f[128] && !f[571]; // c6t596i59
	assign leaf[785] = !f[601] && !f[164] && f[128] && f[571]; // c6t596i59
	assign leaf[786] = !f[601] && f[164]; // c6t596i59
	assign leaf[787] = f[601] && !f[129] && !f[238] && !f[627]; // c6t596i59
	assign leaf[788] = f[601] && !f[129] && !f[238] && f[627]; // c6t596i59
	assign leaf[789] = f[601] && !f[129] && f[238] && !f[99]; // c6t596i59
	assign leaf[790] = f[601] && !f[129] && f[238] && f[99]; // c6t596i59
	assign leaf[791] = f[601] && f[129] && !f[574] && !f[183]; // c6t596i59
	assign leaf[792] = f[601] && f[129] && !f[574] && f[183]; // c6t596i59
	assign leaf[793] = f[601] && f[129] && f[574] && !f[266]; // c6t596i59
	assign leaf[794] = f[601] && f[129] && f[574] && f[266]; // c6t596i59
	assign leaf[795] = !f[205] && !f[467] && !f[326] && !f[123]; // c6t606i60
	assign leaf[796] = !f[205] && !f[467] && !f[326] && f[123]; // c6t606i60
	assign leaf[797] = !f[205] && !f[467] && f[326] && !f[469]; // c6t606i60
	assign leaf[798] = !f[205] && !f[467] && f[326] && f[469]; // c6t606i60
	assign leaf[799] = !f[205] && f[467] && !f[432] && !f[436]; // c6t606i60
	assign leaf[800] = !f[205] && f[467] && !f[432] && f[436]; // c6t606i60
	assign leaf[801] = !f[205] && f[467] && f[432] && !f[287]; // c6t606i60
	assign leaf[802] = !f[205] && f[467] && f[432] && f[287]; // c6t606i60
	assign leaf[803] = f[205] && !f[348] && !f[183] && !f[294]; // c6t606i60
	assign leaf[804] = f[205] && !f[348] && !f[183] && f[294]; // c6t606i60
	assign leaf[805] = f[205] && !f[348] && f[183] && !f[573]; // c6t606i60
	assign leaf[806] = f[205] && !f[348] && f[183] && f[573]; // c6t606i60
	assign leaf[807] = f[205] && f[348] && !f[344] && !f[325]; // c6t606i60
	assign leaf[808] = f[205] && f[348] && !f[344] && f[325]; // c6t606i60
	assign leaf[809] = f[205] && f[348] && f[344] && !f[488]; // c6t606i60
	assign leaf[810] = f[205] && f[348] && f[344] && f[488]; // c6t606i60
	assign leaf[811] = !f[541] && !f[516] && !f[511] && !f[514]; // c6t616i61
	assign leaf[812] = !f[541] && !f[516] && !f[511] && f[514]; // c6t616i61
	assign leaf[813] = !f[541] && !f[516] && f[511] && !f[600]; // c6t616i61
	assign leaf[814] = !f[541] && !f[516] && f[511] && f[600]; // c6t616i61
	assign leaf[815] = !f[541] && f[516] && !f[575] && !f[571]; // c6t616i61
	assign leaf[816] = !f[541] && f[516] && !f[575] && f[571]; // c6t616i61
	assign leaf[817] = !f[541] && f[516] && f[575] && !f[485]; // c6t616i61
	assign leaf[818] = !f[541] && f[516] && f[575] && f[485]; // c6t616i61
	assign leaf[819] = f[541] && !f[401] && !f[291] && !f[237]; // c6t616i61
	assign leaf[820] = f[541] && !f[401] && !f[291] && f[237]; // c6t616i61
	assign leaf[821] = f[541] && !f[401] && f[291] && !f[371]; // c6t616i61
	assign leaf[822] = f[541] && !f[401] && f[291] && f[371]; // c6t616i61
	assign leaf[823] = f[541] && f[401] && !f[457] && !f[403]; // c6t616i61
	assign leaf[824] = f[541] && f[401] && !f[457] && f[403]; // c6t616i61
	assign leaf[825] = f[541] && f[401] && f[457] && !f[136]; // c6t616i61
	assign leaf[826] = f[541] && f[401] && f[457] && f[136]; // c6t616i61
	assign leaf[827] = !f[297] && !f[656] && !f[217] && !f[350]; // c6t626i62
	assign leaf[828] = !f[297] && !f[656] && !f[217] && f[350]; // c6t626i62
	assign leaf[829] = !f[297] && !f[656] && f[217] && !f[580]; // c6t626i62
	assign leaf[830] = !f[297] && !f[656] && f[217] && f[580]; // c6t626i62
	assign leaf[831] = !f[297] && f[656] && !f[355] && !f[152]; // c6t626i62
	assign leaf[832] = !f[297] && f[656] && !f[355] && f[152]; // c6t626i62
	assign leaf[833] = !f[297] && f[656] && f[355] && !f[125]; // c6t626i62
	assign leaf[834] = !f[297] && f[656] && f[355] && f[125]; // c6t626i62
	assign leaf[835] = f[297] && !f[573] && !f[359] && !f[287]; // c6t626i62
	assign leaf[836] = f[297] && !f[573] && !f[359] && f[287]; // c6t626i62
	assign leaf[837] = f[297] && !f[573] && f[359]; // c6t626i62
	assign leaf[838] = f[297] && f[573] && !f[350] && !f[273]; // c6t626i62
	assign leaf[839] = f[297] && f[573] && !f[350] && f[273]; // c6t626i62
	assign leaf[840] = f[297] && f[573] && f[350] && !f[212]; // c6t626i62
	assign leaf[841] = f[297] && f[573] && f[350] && f[212]; // c6t626i62
	assign leaf[842] = !f[268] && !f[349] && !f[686] && !f[322]; // c6t636i63
	assign leaf[843] = !f[268] && !f[349] && !f[686] && f[322]; // c6t636i63
	assign leaf[844] = !f[268] && !f[349] && f[686] && !f[546]; // c6t636i63
	assign leaf[845] = !f[268] && !f[349] && f[686] && f[546]; // c6t636i63
	assign leaf[846] = !f[268] && f[349] && !f[123] && !f[629]; // c6t636i63
	assign leaf[847] = !f[268] && f[349] && !f[123] && f[629]; // c6t636i63
	assign leaf[848] = !f[268] && f[349] && f[123] && !f[599]; // c6t636i63
	assign leaf[849] = !f[268] && f[349] && f[123] && f[599]; // c6t636i63
	assign leaf[850] = f[268] && !f[408] && !f[570] && !f[239]; // c6t636i63
	assign leaf[851] = f[268] && !f[408] && !f[570] && f[239]; // c6t636i63
	assign leaf[852] = f[268] && !f[408] && f[570] && !f[490]; // c6t636i63
	assign leaf[853] = f[268] && !f[408] && f[570] && f[490]; // c6t636i63
	assign leaf[854] = f[268] && f[408] && !f[349] && !f[606]; // c6t636i63
	assign leaf[855] = f[268] && f[408] && !f[349] && f[606]; // c6t636i63
	assign leaf[856] = f[268] && f[408] && f[349] && !f[579]; // c6t636i63
	assign leaf[857] = f[268] && f[408] && f[349] && f[579]; // c6t636i63
	assign leaf[858] = !f[101] && !f[275] && !f[205] && !f[467]; // c6t646i64
	assign leaf[859] = !f[101] && !f[275] && !f[205] && f[467]; // c6t646i64
	assign leaf[860] = !f[101] && !f[275] && f[205] && !f[182]; // c6t646i64
	assign leaf[861] = !f[101] && !f[275] && f[205] && f[182]; // c6t646i64
	assign leaf[862] = !f[101] && f[275] && !f[605]; // c6t646i64
	assign leaf[863] = !f[101] && f[275] && f[605]; // c6t646i64
	assign leaf[864] = f[101] && !f[127] && !f[570]; // c6t646i64
	assign leaf[865] = f[101] && !f[127] && f[570] && !f[238]; // c6t646i64
	assign leaf[866] = f[101] && !f[127] && f[570] && f[238]; // c6t646i64
	assign leaf[867] = f[101] && f[127] && !f[547] && !f[605]; // c6t646i64
	assign leaf[868] = f[101] && f[127] && !f[547] && f[605]; // c6t646i64
	assign leaf[869] = f[101] && f[127] && f[547] && !f[539]; // c6t646i64
	assign leaf[870] = f[101] && f[127] && f[547] && f[539]; // c6t646i64
	assign leaf[871] = !f[268] && !f[136] && !f[231] && !f[636]; // c6t656i65
	assign leaf[872] = !f[268] && !f[136] && !f[231] && f[636]; // c6t656i65
	assign leaf[873] = !f[268] && !f[136] && f[231] && !f[347]; // c6t656i65
	assign leaf[874] = !f[268] && !f[136] && f[231] && f[347]; // c6t656i65
	assign leaf[875] = !f[268] && f[136]; // c6t656i65
	assign leaf[876] = f[268] && !f[380] && !f[570] && !f[512]; // c6t656i65
	assign leaf[877] = f[268] && !f[380] && !f[570] && f[512]; // c6t656i65
	assign leaf[878] = f[268] && !f[380] && f[570] && !f[490]; // c6t656i65
	assign leaf[879] = f[268] && !f[380] && f[570] && f[490]; // c6t656i65
	assign leaf[880] = f[268] && f[380] && !f[324] && !f[486]; // c6t656i65
	assign leaf[881] = f[268] && f[380] && !f[324] && f[486]; // c6t656i65
	assign leaf[882] = f[268] && f[380] && f[324] && !f[161]; // c6t656i65
	assign leaf[883] = f[268] && f[380] && f[324] && f[161]; // c6t656i65
	assign leaf[884] = !f[91] && !f[213] && !f[324] && !f[323]; // c6t666i66
	assign leaf[885] = !f[91] && !f[213] && !f[324] && f[323]; // c6t666i66
	assign leaf[886] = !f[91] && !f[213] && f[324] && !f[238]; // c6t666i66
	assign leaf[887] = !f[91] && !f[213] && f[324] && f[238]; // c6t666i66
	assign leaf[888] = !f[91] && f[213] && !f[325] && !f[356]; // c6t666i66
	assign leaf[889] = !f[91] && f[213] && !f[325] && f[356]; // c6t666i66
	assign leaf[890] = !f[91] && f[213] && f[325] && !f[190]; // c6t666i66
	assign leaf[891] = !f[91] && f[213] && f[325] && f[190]; // c6t666i66
	assign leaf[892] = f[91]; // c6t666i66
	assign leaf[893] = !f[602] && !f[126] && !f[629] && !f[291]; // c6t676i67
	assign leaf[894] = !f[602] && !f[126] && !f[629] && f[291]; // c6t676i67
	assign leaf[895] = !f[602] && !f[126] && f[629] && !f[522]; // c6t676i67
	assign leaf[896] = !f[602] && !f[126] && f[629] && f[522]; // c6t676i67
	assign leaf[897] = !f[602] && f[126] && !f[574] && !f[491]; // c6t676i67
	assign leaf[898] = !f[602] && f[126] && !f[574] && f[491]; // c6t676i67
	assign leaf[899] = !f[602] && f[126] && f[574] && !f[208]; // c6t676i67
	assign leaf[900] = !f[602] && f[126] && f[574] && f[208]; // c6t676i67
	assign leaf[901] = f[602] && !f[486] && !f[543] && !f[544]; // c6t676i67
	assign leaf[902] = f[602] && !f[486] && !f[543] && f[544]; // c6t676i67
	assign leaf[903] = f[602] && !f[486] && f[543] && !f[426]; // c6t676i67
	assign leaf[904] = f[602] && !f[486] && f[543] && f[426]; // c6t676i67
	assign leaf[905] = f[602] && f[486] && !f[189] && !f[374]; // c6t676i67
	assign leaf[906] = f[602] && f[486] && !f[189] && f[374]; // c6t676i67
	assign leaf[907] = f[602] && f[486] && f[189] && !f[521]; // c6t676i67
	assign leaf[908] = f[602] && f[486] && f[189] && f[521]; // c6t676i67
	assign leaf[909] = !f[270] && !f[514] && !f[406] && !f[267]; // c6t686i68
	assign leaf[910] = !f[270] && !f[514] && !f[406] && f[267]; // c6t686i68
	assign leaf[911] = !f[270] && !f[514] && f[406] && !f[462]; // c6t686i68
	assign leaf[912] = !f[270] && !f[514] && f[406] && f[462]; // c6t686i68
	assign leaf[913] = !f[270] && f[514] && !f[401] && !f[153]; // c6t686i68
	assign leaf[914] = !f[270] && f[514] && !f[401] && f[153]; // c6t686i68
	assign leaf[915] = !f[270] && f[514] && f[401] && !f[571]; // c6t686i68
	assign leaf[916] = !f[270] && f[514] && f[401] && f[571]; // c6t686i68
	assign leaf[917] = f[270] && !f[272] && !f[541] && !f[325]; // c6t686i68
	assign leaf[918] = f[270] && !f[272] && !f[541] && f[325]; // c6t686i68
	assign leaf[919] = f[270] && !f[272] && f[541] && !f[540]; // c6t686i68
	assign leaf[920] = f[270] && !f[272] && f[541] && f[540]; // c6t686i68
	assign leaf[921] = f[270] && f[272] && !f[186] && !f[355]; // c6t686i68
	assign leaf[922] = f[270] && f[272] && !f[186] && f[355]; // c6t686i68
	assign leaf[923] = f[270] && f[272] && f[186] && !f[468]; // c6t686i68
	assign leaf[924] = f[270] && f[272] && f[186] && f[468]; // c6t686i68
	assign leaf[925] = !f[601] && !f[208] && !f[523] && !f[542]; // c6t696i69
	assign leaf[926] = !f[601] && !f[208] && !f[523] && f[542]; // c6t696i69
	assign leaf[927] = !f[601] && !f[208] && f[523] && !f[263]; // c6t696i69
	assign leaf[928] = !f[601] && !f[208] && f[523] && f[263]; // c6t696i69
	assign leaf[929] = !f[601] && f[208] && !f[180]; // c6t696i69
	assign leaf[930] = !f[601] && f[208] && f[180] && !f[263]; // c6t696i69
	assign leaf[931] = !f[601] && f[208] && f[180] && f[263]; // c6t696i69
	assign leaf[932] = f[601] && !f[627] && !f[178] && !f[516]; // c6t696i69
	assign leaf[933] = f[601] && !f[627] && !f[178] && f[516]; // c6t696i69
	assign leaf[934] = f[601] && !f[627] && f[178] && !f[631]; // c6t696i69
	assign leaf[935] = f[601] && !f[627] && f[178] && f[631]; // c6t696i69
	assign leaf[936] = f[601] && f[627] && !f[127] && !f[209]; // c6t696i69
	assign leaf[937] = f[601] && f[627] && !f[127] && f[209]; // c6t696i69
	assign leaf[938] = f[601] && f[627] && f[127] && !f[455]; // c6t696i69
	assign leaf[939] = f[601] && f[627] && f[127] && f[455]; // c6t696i69
	assign leaf[940] = !f[236] && !f[181] && !f[656] && !f[480]; // c6t706i70
	assign leaf[941] = !f[236] && !f[181] && !f[656] && f[480]; // c6t706i70
	assign leaf[942] = !f[236] && !f[181] && f[656] && !f[547]; // c6t706i70
	assign leaf[943] = !f[236] && !f[181] && f[656] && f[547]; // c6t706i70
	assign leaf[944] = !f[236] && f[181] && !f[516] && !f[357]; // c6t706i70
	assign leaf[945] = !f[236] && f[181] && !f[516] && f[357]; // c6t706i70
	assign leaf[946] = !f[236] && f[181] && f[516] && !f[184]; // c6t706i70
	assign leaf[947] = !f[236] && f[181] && f[516] && f[184]; // c6t706i70
	assign leaf[948] = f[236] && !f[541] && !f[347] && !f[539]; // c6t706i70
	assign leaf[949] = f[236] && !f[541] && !f[347] && f[539]; // c6t706i70
	assign leaf[950] = f[236] && !f[541] && f[347] && !f[487]; // c6t706i70
	assign leaf[951] = f[236] && !f[541] && f[347] && f[487]; // c6t706i70
	assign leaf[952] = f[236] && f[541] && !f[401] && !f[371]; // c6t706i70
	assign leaf[953] = f[236] && f[541] && !f[401] && f[371]; // c6t706i70
	assign leaf[954] = f[236] && f[541] && f[401] && !f[128]; // c6t706i70
	assign leaf[955] = f[236] && f[541] && f[401] && f[128]; // c6t706i70
	assign leaf[956] = !f[622] && !f[101] && !f[212] && !f[320]; // c6t716i71
	assign leaf[957] = !f[622] && !f[101] && !f[212] && f[320]; // c6t716i71
	assign leaf[958] = !f[622] && !f[101] && f[212] && !f[486]; // c6t716i71
	assign leaf[959] = !f[622] && !f[101] && f[212] && f[486]; // c6t716i71
	assign leaf[960] = !f[622] && f[101] && !f[211] && !f[580]; // c6t716i71
	assign leaf[961] = !f[622] && f[101] && !f[211] && f[580]; // c6t716i71
	assign leaf[962] = !f[622] && f[101] && f[211] && !f[631]; // c6t716i71
	assign leaf[963] = !f[622] && f[101] && f[211] && f[631]; // c6t716i71
	assign leaf[964] = f[622]; // c6t716i71
	assign leaf[965] = !f[269] && !f[301] && !f[232] && !f[399]; // c6t726i72
	assign leaf[966] = !f[269] && !f[301] && !f[232] && f[399]; // c6t726i72
	assign leaf[967] = !f[269] && !f[301] && f[232] && !f[347]; // c6t726i72
	assign leaf[968] = !f[269] && !f[301] && f[232] && f[347]; // c6t726i72
	assign leaf[969] = !f[269] && f[301] && !f[299] && !f[359]; // c6t726i72
	assign leaf[970] = !f[269] && f[301] && !f[299] && f[359]; // c6t726i72
	assign leaf[971] = !f[269] && f[301] && f[299] && !f[383]; // c6t726i72
	assign leaf[972] = !f[269] && f[301] && f[299] && f[383]; // c6t726i72
	assign leaf[973] = f[269] && !f[662] && !f[164] && !f[604]; // c6t726i72
	assign leaf[974] = f[269] && !f[662] && !f[164] && f[604]; // c6t726i72
	assign leaf[975] = f[269] && !f[662] && f[164] && !f[319]; // c6t726i72
	assign leaf[976] = f[269] && !f[662] && f[164] && f[319]; // c6t726i72
	assign leaf[977] = f[269] && f[662]; // c6t726i72
	assign leaf[978] = !f[432] && !f[214] && !f[349] && !f[155]; // c6t736i73
	assign leaf[979] = !f[432] && !f[214] && !f[349] && f[155]; // c6t736i73
	assign leaf[980] = !f[432] && !f[214] && f[349] && !f[457]; // c6t736i73
	assign leaf[981] = !f[432] && !f[214] && f[349] && f[457]; // c6t736i73
	assign leaf[982] = !f[432] && f[214] && !f[238] && !f[433]; // c6t736i73
	assign leaf[983] = !f[432] && f[214] && !f[238] && f[433]; // c6t736i73
	assign leaf[984] = !f[432] && f[214] && f[238] && !f[159]; // c6t736i73
	assign leaf[985] = !f[432] && f[214] && f[238] && f[159]; // c6t736i73
	assign leaf[986] = f[432] && !f[516] && !f[541] && !f[510]; // c6t736i73
	assign leaf[987] = f[432] && !f[516] && !f[541] && f[510]; // c6t736i73
	assign leaf[988] = f[432] && !f[516] && f[541] && !f[326]; // c6t736i73
	assign leaf[989] = f[432] && !f[516] && f[541] && f[326]; // c6t736i73
	assign leaf[990] = f[432] && f[516] && !f[155] && !f[237]; // c6t736i73
	assign leaf[991] = f[432] && f[516] && !f[155] && f[237]; // c6t736i73
	assign leaf[992] = f[432] && f[516] && f[155] && !f[244]; // c6t736i73
	assign leaf[993] = f[432] && f[516] && f[155] && f[244]; // c6t736i73
	assign leaf[994] = !f[302] && !f[299] && !f[399] && !f[518]; // c6t746i74
	assign leaf[995] = !f[302] && !f[299] && !f[399] && f[518]; // c6t746i74
	assign leaf[996] = !f[302] && !f[299] && f[399] && !f[269]; // c6t746i74
	assign leaf[997] = !f[302] && !f[299] && f[399] && f[269]; // c6t746i74
	assign leaf[998] = !f[302] && f[299] && !f[457] && !f[301]; // c6t746i74
	assign leaf[999] = !f[302] && f[299] && !f[457] && f[301]; // c6t746i74
	assign leaf[1000] = !f[302] && f[299] && f[457] && !f[382]; // c6t746i74
	assign leaf[1001] = !f[302] && f[299] && f[457] && f[382]; // c6t746i74
	assign leaf[1002] = f[302] && !f[416] && !f[271] && !f[408]; // c6t746i74
	assign leaf[1003] = f[302] && !f[416] && !f[271] && f[408]; // c6t746i74
	assign leaf[1004] = f[302] && !f[416] && f[271] && !f[430]; // c6t746i74
	assign leaf[1005] = f[302] && !f[416] && f[271] && f[430]; // c6t746i74
	assign leaf[1006] = f[302] && f[416]; // c6t746i74
	assign leaf[1007] = !f[652] && !f[655] && !f[162] && !f[374]; // c6t756i75
	assign leaf[1008] = !f[652] && !f[655] && !f[162] && f[374]; // c6t756i75
	assign leaf[1009] = !f[652] && !f[655] && f[162] && !f[189]; // c6t756i75
	assign leaf[1010] = !f[652] && !f[655] && f[162] && f[189]; // c6t756i75
	assign leaf[1011] = !f[652] && f[655] && !f[241] && !f[211]; // c6t756i75
	assign leaf[1012] = !f[652] && f[655] && !f[241] && f[211]; // c6t756i75
	assign leaf[1013] = !f[652] && f[655] && f[241] && !f[379]; // c6t756i75
	assign leaf[1014] = !f[652] && f[655] && f[241] && f[379]; // c6t756i75
	assign leaf[1015] = f[652] && !f[488]; // c6t756i75
	assign leaf[1016] = f[652] && f[488]; // c6t756i75
	assign leaf[1017] = !f[682] && !f[638] && !f[610] && !f[406]; // c6t766i76
	assign leaf[1018] = !f[682] && !f[638] && !f[610] && f[406]; // c6t766i76
	assign leaf[1019] = !f[682] && !f[638] && f[610] && !f[315]; // c6t766i76
	assign leaf[1020] = !f[682] && !f[638] && f[610] && f[315]; // c6t766i76
	assign leaf[1021] = !f[682] && f[638]; // c6t766i76
	assign leaf[1022] = f[682]; // c6t766i76
	assign leaf[1023] = !f[214] && !f[637] && !f[295] && !f[247]; // c6t776i77
	assign leaf[1024] = !f[214] && !f[637] && !f[295] && f[247]; // c6t776i77
	assign leaf[1025] = !f[214] && !f[637] && f[295] && !f[265]; // c6t776i77
	assign leaf[1026] = !f[214] && !f[637] && f[295] && f[265]; // c6t776i77
	assign leaf[1027] = !f[214] && f[637]; // c6t776i77
	assign leaf[1028] = f[214] && !f[348] && !f[377] && !f[320]; // c6t776i77
	assign leaf[1029] = f[214] && !f[348] && !f[377] && f[320]; // c6t776i77
	assign leaf[1030] = f[214] && !f[348] && f[377] && !f[316]; // c6t776i77
	assign leaf[1031] = f[214] && !f[348] && f[377] && f[316]; // c6t776i77
	assign leaf[1032] = f[214] && f[348] && !f[687] && !f[235]; // c6t776i77
	assign leaf[1033] = f[214] && f[348] && !f[687] && f[235]; // c6t776i77
	assign leaf[1034] = f[214] && f[348] && f[687]; // c6t776i77
	assign leaf[1035] = !f[571] && !f[574] && !f[541] && !f[578]; // c6t786i78
	assign leaf[1036] = !f[571] && !f[574] && !f[541] && f[578]; // c6t786i78
	assign leaf[1037] = !f[571] && !f[574] && f[541] && !f[384]; // c6t786i78
	assign leaf[1038] = !f[571] && !f[574] && f[541] && f[384]; // c6t786i78
	assign leaf[1039] = !f[571] && f[574] && !f[156] && !f[270]; // c6t786i78
	assign leaf[1040] = !f[571] && f[574] && !f[156] && f[270]; // c6t786i78
	assign leaf[1041] = !f[571] && f[574] && f[156] && !f[100]; // c6t786i78
	assign leaf[1042] = !f[571] && f[574] && f[156] && f[100]; // c6t786i78
	assign leaf[1043] = f[571] && !f[486] && !f[426] && !f[262]; // c6t786i78
	assign leaf[1044] = f[571] && !f[486] && !f[426] && f[262]; // c6t786i78
	assign leaf[1045] = f[571] && !f[486] && f[426] && !f[272]; // c6t786i78
	assign leaf[1046] = f[571] && !f[486] && f[426] && f[272]; // c6t786i78
	assign leaf[1047] = f[571] && f[486] && !f[540] && !f[514]; // c6t786i78
	assign leaf[1048] = f[571] && f[486] && !f[540] && f[514]; // c6t786i78
	assign leaf[1049] = f[571] && f[486] && f[540] && !f[400]; // c6t786i78
	assign leaf[1050] = f[571] && f[486] && f[540] && f[400]; // c6t786i78
	assign leaf[1051] = !f[445] && !f[234] && !f[151] && !f[96]; // c6t796i79
	assign leaf[1052] = !f[445] && !f[234] && !f[151] && f[96]; // c6t796i79
	assign leaf[1053] = !f[445] && !f[234] && f[151] && !f[518]; // c6t796i79
	assign leaf[1054] = !f[445] && !f[234] && f[151] && f[518]; // c6t796i79
	assign leaf[1055] = !f[445] && f[234] && !f[373] && !f[426]; // c6t796i79
	assign leaf[1056] = !f[445] && f[234] && !f[373] && f[426]; // c6t796i79
	assign leaf[1057] = !f[445] && f[234] && f[373] && !f[152]; // c6t796i79
	assign leaf[1058] = !f[445] && f[234] && f[373] && f[152]; // c6t796i79
	assign leaf[1059] = f[445]; // c6t796i79
	assign leaf[1060] = !f[517] && !f[234] && !f[151] && !f[242]; // c6t806i80
	assign leaf[1061] = !f[517] && !f[234] && !f[151] && f[242]; // c6t806i80
	assign leaf[1062] = !f[517] && !f[234] && f[151] && !f[347]; // c6t806i80
	assign leaf[1063] = !f[517] && !f[234] && f[151] && f[347]; // c6t806i80
	assign leaf[1064] = !f[517] && f[234] && !f[428] && !f[436]; // c6t806i80
	assign leaf[1065] = !f[517] && f[234] && !f[428] && f[436]; // c6t806i80
	assign leaf[1066] = !f[517] && f[234] && f[428] && !f[601]; // c6t806i80
	assign leaf[1067] = !f[517] && f[234] && f[428] && f[601]; // c6t806i80
	assign leaf[1068] = f[517] && !f[212] && !f[246] && !f[383]; // c6t806i80
	assign leaf[1069] = f[517] && !f[212] && !f[246] && f[383]; // c6t806i80
	assign leaf[1070] = f[517] && !f[212] && f[246] && !f[406]; // c6t806i80
	assign leaf[1071] = f[517] && !f[212] && f[246] && f[406]; // c6t806i80
	assign leaf[1072] = f[517] && f[212] && !f[599] && !f[551]; // c6t806i80
	assign leaf[1073] = f[517] && f[212] && !f[599] && f[551]; // c6t806i80
	assign leaf[1074] = f[517] && f[212] && f[599] && !f[521]; // c6t806i80
	assign leaf[1075] = f[517] && f[212] && f[599] && f[521]; // c6t806i80
	assign leaf[1076] = !f[459] && !f[515] && !f[489] && !f[512]; // c6t816i81
	assign leaf[1077] = !f[459] && !f[515] && !f[489] && f[512]; // c6t816i81
	assign leaf[1078] = !f[459] && !f[515] && f[489] && !f[405]; // c6t816i81
	assign leaf[1079] = !f[459] && !f[515] && f[489] && f[405]; // c6t816i81
	assign leaf[1080] = !f[459] && f[515] && !f[359] && !f[457]; // c6t816i81
	assign leaf[1081] = !f[459] && f[515] && !f[359] && f[457]; // c6t816i81
	assign leaf[1082] = !f[459] && f[515] && f[359] && !f[407]; // c6t816i81
	assign leaf[1083] = !f[459] && f[515] && f[359] && f[407]; // c6t816i81
	assign leaf[1084] = f[459] && !f[610] && !f[316] && !f[687]; // c6t816i81
	assign leaf[1085] = f[459] && !f[610] && !f[316] && f[687]; // c6t816i81
	assign leaf[1086] = f[459] && !f[610] && f[316] && !f[384]; // c6t816i81
	assign leaf[1087] = f[459] && !f[610] && f[316] && f[384]; // c6t816i81
	assign leaf[1088] = f[459] && f[610]; // c6t816i81
	assign leaf[1089] = !f[652] && !f[267] && !f[237] && !f[183]; // c6t826i82
	assign leaf[1090] = !f[652] && !f[267] && !f[237] && f[183]; // c6t826i82
	assign leaf[1091] = !f[652] && !f[267] && f[237] && !f[328]; // c6t826i82
	assign leaf[1092] = !f[652] && !f[267] && f[237] && f[328]; // c6t826i82
	assign leaf[1093] = !f[652] && f[267] && !f[321] && !f[545]; // c6t826i82
	assign leaf[1094] = !f[652] && f[267] && !f[321] && f[545]; // c6t826i82
	assign leaf[1095] = !f[652] && f[267] && f[321] && !f[580]; // c6t826i82
	assign leaf[1096] = !f[652] && f[267] && f[321] && f[580]; // c6t826i82
	assign leaf[1097] = f[652] && !f[512]; // c6t826i82
	assign leaf[1098] = f[652] && f[512]; // c6t826i82
	assign leaf[1099] = !f[299] && !f[301] && !f[272] && !f[383]; // c6t836i83
	assign leaf[1100] = !f[299] && !f[301] && !f[272] && f[383]; // c6t836i83
	assign leaf[1101] = !f[299] && !f[301] && f[272]; // c6t836i83
	assign leaf[1102] = !f[299] && f[301] && !f[403] && !f[434]; // c6t836i83
	assign leaf[1103] = !f[299] && f[301] && !f[403] && f[434]; // c6t836i83
	assign leaf[1104] = !f[299] && f[301] && f[403]; // c6t836i83
	assign leaf[1105] = f[299] && !f[382] && !f[658] && !f[388]; // c6t836i83
	assign leaf[1106] = f[299] && !f[382] && !f[658] && f[388]; // c6t836i83
	assign leaf[1107] = f[299] && !f[382] && f[658] && !f[293]; // c6t836i83
	assign leaf[1108] = f[299] && !f[382] && f[658] && f[293]; // c6t836i83
	assign leaf[1109] = f[299] && f[382] && !f[352] && !f[301]; // c6t836i83
	assign leaf[1110] = f[299] && f[382] && !f[352] && f[301]; // c6t836i83
	assign leaf[1111] = f[299] && f[382] && f[352] && !f[494]; // c6t836i83
	assign leaf[1112] = f[299] && f[382] && f[352] && f[494]; // c6t836i83
	assign leaf[1113] = !f[571] && !f[575] && !f[399] && !f[187]; // c6t846i84
	assign leaf[1114] = !f[571] && !f[575] && !f[399] && f[187]; // c6t846i84
	assign leaf[1115] = !f[571] && !f[575] && f[399] && !f[401]; // c6t846i84
	assign leaf[1116] = !f[571] && !f[575] && f[399] && f[401]; // c6t846i84
	assign leaf[1117] = !f[571] && f[575] && !f[659] && !f[242]; // c6t846i84
	assign leaf[1118] = !f[571] && f[575] && !f[659] && f[242]; // c6t846i84
	assign leaf[1119] = !f[571] && f[575] && f[659] && !f[545]; // c6t846i84
	assign leaf[1120] = !f[571] && f[575] && f[659] && f[545]; // c6t846i84
	assign leaf[1121] = f[571] && !f[486] && !f[181] && !f[98]; // c6t846i84
	assign leaf[1122] = f[571] && !f[486] && !f[181] && f[98]; // c6t846i84
	assign leaf[1123] = f[571] && !f[486] && f[181] && !f[315]; // c6t846i84
	assign leaf[1124] = f[571] && !f[486] && f[181] && f[315]; // c6t846i84
	assign leaf[1125] = f[571] && f[486] && !f[687] && !f[568]; // c6t846i84
	assign leaf[1126] = f[571] && f[486] && !f[687] && f[568]; // c6t846i84
	assign leaf[1127] = f[571] && f[486] && f[687]; // c6t846i84
	assign leaf[1128] = !f[247] && !f[574] && !f[570] && !f[571]; // c6t856i85
	assign leaf[1129] = !f[247] && !f[574] && !f[570] && f[571]; // c6t856i85
	assign leaf[1130] = !f[247] && !f[574] && f[570] && !f[152]; // c6t856i85
	assign leaf[1131] = !f[247] && !f[574] && f[570] && f[152]; // c6t856i85
	assign leaf[1132] = !f[247] && f[574] && !f[209] && !f[320]; // c6t856i85
	assign leaf[1133] = !f[247] && f[574] && !f[209] && f[320]; // c6t856i85
	assign leaf[1134] = !f[247] && f[574] && f[209] && !f[126]; // c6t856i85
	assign leaf[1135] = !f[247] && f[574] && f[209] && f[126]; // c6t856i85
	assign leaf[1136] = f[247] && !f[630]; // c6t856i85
	assign leaf[1137] = f[247] && f[630]; // c6t856i85
	assign leaf[1138] = !f[107] && !f[214] && !f[293] && !f[155]; // c6t866i86
	assign leaf[1139] = !f[107] && !f[214] && !f[293] && f[155]; // c6t866i86
	assign leaf[1140] = !f[107] && !f[214] && f[293] && !f[156]; // c6t866i86
	assign leaf[1141] = !f[107] && !f[214] && f[293] && f[156]; // c6t866i86
	assign leaf[1142] = !f[107] && f[214] && !f[433] && !f[509]; // c6t866i86
	assign leaf[1143] = !f[107] && f[214] && !f[433] && f[509]; // c6t866i86
	assign leaf[1144] = !f[107] && f[214] && f[433] && !f[352]; // c6t866i86
	assign leaf[1145] = !f[107] && f[214] && f[433] && f[352]; // c6t866i86
	assign leaf[1146] = f[107]; // c6t866i86
	assign leaf[1147] = !f[299] && !f[301] && !f[383] && !f[123]; // c6t876i87
	assign leaf[1148] = !f[299] && !f[301] && !f[383] && f[123]; // c6t876i87
	assign leaf[1149] = !f[299] && !f[301] && f[383] && !f[405]; // c6t876i87
	assign leaf[1150] = !f[299] && !f[301] && f[383] && f[405]; // c6t876i87
	assign leaf[1151] = !f[299] && f[301] && !f[489]; // c6t876i87
	assign leaf[1152] = !f[299] && f[301] && f[489] && !f[289]; // c6t876i87
	assign leaf[1153] = !f[299] && f[301] && f[489] && f[289]; // c6t876i87
	assign leaf[1154] = f[299] && !f[358] && !f[348] && !f[233]; // c6t876i87
	assign leaf[1155] = f[299] && !f[358] && !f[348] && f[233]; // c6t876i87
	assign leaf[1156] = f[299] && !f[358] && f[348] && !f[542]; // c6t876i87
	assign leaf[1157] = f[299] && !f[358] && f[348] && f[542]; // c6t876i87
	assign leaf[1158] = f[299] && f[358] && !f[600]; // c6t876i87
	assign leaf[1159] = f[299] && f[358] && f[600] && !f[486]; // c6t876i87
	assign leaf[1160] = f[299] && f[358] && f[600] && f[486]; // c6t876i87
	assign leaf[1161] = !f[629] && !f[383] && !f[549] && !f[521]; // c6t886i88
	assign leaf[1162] = !f[629] && !f[383] && !f[549] && f[521]; // c6t886i88
	assign leaf[1163] = !f[629] && !f[383] && f[549] && !f[514]; // c6t886i88
	assign leaf[1164] = !f[629] && !f[383] && f[549] && f[514]; // c6t886i88
	assign leaf[1165] = !f[629] && f[383] && !f[273] && !f[547]; // c6t886i88
	assign leaf[1166] = !f[629] && f[383] && !f[273] && f[547]; // c6t886i88
	assign leaf[1167] = !f[629] && f[383] && f[273]; // c6t886i88
	assign leaf[1168] = f[629] && !f[260] && !f[608] && !f[687]; // c6t886i88
	assign leaf[1169] = f[629] && !f[260] && !f[608] && f[687]; // c6t886i88
	assign leaf[1170] = f[629] && !f[260] && f[608] && !f[428]; // c6t886i88
	assign leaf[1171] = f[629] && !f[260] && f[608] && f[428]; // c6t886i88
	assign leaf[1172] = f[629] && f[260] && !f[464] && !f[545]; // c6t886i88
	assign leaf[1173] = f[629] && f[260] && !f[464] && f[545]; // c6t886i88
	assign leaf[1174] = f[629] && f[260] && f[464] && !f[483]; // c6t886i88
	assign leaf[1175] = f[629] && f[260] && f[464] && f[483]; // c6t886i88
	assign leaf[1176] = !f[409] && !f[436] && !f[354] && !f[603]; // c6t896i89
	assign leaf[1177] = !f[409] && !f[436] && !f[354] && f[603]; // c6t896i89
	assign leaf[1178] = !f[409] && !f[436] && f[354] && !f[270]; // c6t896i89
	assign leaf[1179] = !f[409] && !f[436] && f[354] && f[270]; // c6t896i89
	assign leaf[1180] = !f[409] && f[436] && !f[576] && !f[440]; // c6t896i89
	assign leaf[1181] = !f[409] && f[436] && !f[576] && f[440]; // c6t896i89
	assign leaf[1182] = !f[409] && f[436] && f[576] && !f[406]; // c6t896i89
	assign leaf[1183] = !f[409] && f[436] && f[576] && f[406]; // c6t896i89
	assign leaf[1184] = f[409] && !f[435] && !f[326] && !f[429]; // c6t896i89
	assign leaf[1185] = f[409] && !f[435] && !f[326] && f[429]; // c6t896i89
	assign leaf[1186] = f[409] && !f[435] && f[326] && !f[239]; // c6t896i89
	assign leaf[1187] = f[409] && !f[435] && f[326] && f[239]; // c6t896i89
	assign leaf[1188] = f[409] && f[435] && !f[627] && !f[545]; // c6t896i89
	assign leaf[1189] = f[409] && f[435] && !f[627] && f[545]; // c6t896i89
	assign leaf[1190] = f[409] && f[435] && f[627] && !f[464]; // c6t896i89
	assign leaf[1191] = f[409] && f[435] && f[627] && f[464]; // c6t896i89
	assign leaf[1192] = !f[355] && !f[272] && !f[297] && !f[358]; // c6t906i90
	assign leaf[1193] = !f[355] && !f[272] && !f[297] && f[358]; // c6t906i90
	assign leaf[1194] = !f[355] && !f[272] && f[297] && !f[625]; // c6t906i90
	assign leaf[1195] = !f[355] && !f[272] && f[297] && f[625]; // c6t906i90
	assign leaf[1196] = !f[355] && f[272] && !f[635] && !f[291]; // c6t906i90
	assign leaf[1197] = !f[355] && f[272] && !f[635] && f[291]; // c6t906i90
	assign leaf[1198] = !f[355] && f[272] && f[635]; // c6t906i90
	assign leaf[1199] = f[355] && !f[352] && !f[441] && !f[358]; // c6t906i90
	assign leaf[1200] = f[355] && !f[352] && !f[441] && f[358]; // c6t906i90
	assign leaf[1201] = f[355] && !f[352] && f[441] && !f[456]; // c6t906i90
	assign leaf[1202] = f[355] && !f[352] && f[441] && f[456]; // c6t906i90
	assign leaf[1203] = f[355] && f[352] && !f[349] && !f[239]; // c6t906i90
	assign leaf[1204] = f[355] && f[352] && !f[349] && f[239]; // c6t906i90
	assign leaf[1205] = f[355] && f[352] && f[349] && !f[400]; // c6t906i90
	assign leaf[1206] = f[355] && f[352] && f[349] && f[400]; // c6t906i90
	assign leaf[1207] = !f[516] && !f[485] && !f[483] && !f[486]; // c6t916i91
	assign leaf[1208] = !f[516] && !f[485] && !f[483] && f[486]; // c6t916i91
	assign leaf[1209] = !f[516] && !f[485] && f[483] && !f[497]; // c6t916i91
	assign leaf[1210] = !f[516] && !f[485] && f[483] && f[497]; // c6t916i91
	assign leaf[1211] = !f[516] && f[485] && !f[373] && !f[262]; // c6t916i91
	assign leaf[1212] = !f[516] && f[485] && !f[373] && f[262]; // c6t916i91
	assign leaf[1213] = !f[516] && f[485] && f[373] && !f[241]; // c6t916i91
	assign leaf[1214] = !f[516] && f[485] && f[373] && f[241]; // c6t916i91
	assign leaf[1215] = f[516] && !f[275] && !f[216] && !f[294]; // c6t916i91
	assign leaf[1216] = f[516] && !f[275] && !f[216] && f[294]; // c6t916i91
	assign leaf[1217] = f[516] && !f[275] && f[216] && !f[380]; // c6t916i91
	assign leaf[1218] = f[516] && !f[275] && f[216] && f[380]; // c6t916i91
	assign leaf[1219] = f[516] && f[275]; // c6t916i91
	assign leaf[1220] = !f[522] && !f[570] && !f[634] && !f[242]; // c6t926i92
	assign leaf[1221] = !f[522] && !f[570] && !f[634] && f[242]; // c6t926i92
	assign leaf[1222] = !f[522] && !f[570] && f[634] && !f[184]; // c6t926i92
	assign leaf[1223] = !f[522] && !f[570] && f[634] && f[184]; // c6t926i92
	assign leaf[1224] = !f[522] && f[570] && !f[408] && !f[434]; // c6t926i92
	assign leaf[1225] = !f[522] && f[570] && !f[408] && f[434]; // c6t926i92
	assign leaf[1226] = !f[522] && f[570] && f[408] && !f[466]; // c6t926i92
	assign leaf[1227] = !f[522] && f[570] && f[408] && f[466]; // c6t926i92
	assign leaf[1228] = f[522] && !f[261] && !f[151] && !f[217]; // c6t926i92
	assign leaf[1229] = f[522] && !f[261] && !f[151] && f[217]; // c6t926i92
	assign leaf[1230] = f[522] && !f[261] && f[151] && !f[239]; // c6t926i92
	assign leaf[1231] = f[522] && !f[261] && f[151] && f[239]; // c6t926i92
	assign leaf[1232] = f[522] && f[261] && !f[264] && !f[459]; // c6t926i92
	assign leaf[1233] = f[522] && f[261] && !f[264] && f[459]; // c6t926i92
	assign leaf[1234] = f[522] && f[261] && f[264] && !f[125]; // c6t926i92
	assign leaf[1235] = f[522] && f[261] && f[264] && f[125]; // c6t926i92
	assign leaf[1236] = !f[516] && !f[486] && !f[511] && !f[485]; // c6t936i93
	assign leaf[1237] = !f[516] && !f[486] && !f[511] && f[485]; // c6t936i93
	assign leaf[1238] = !f[516] && !f[486] && f[511] && !f[349]; // c6t936i93
	assign leaf[1239] = !f[516] && !f[486] && f[511] && f[349]; // c6t936i93
	assign leaf[1240] = !f[516] && f[486] && !f[542] && !f[133]; // c6t936i93
	assign leaf[1241] = !f[516] && f[486] && !f[542] && f[133]; // c6t936i93
	assign leaf[1242] = !f[516] && f[486] && f[542] && !f[295]; // c6t936i93
	assign leaf[1243] = !f[516] && f[486] && f[542] && f[295]; // c6t936i93
	assign leaf[1244] = f[516] && !f[432] && !f[515] && !f[380]; // c6t936i93
	assign leaf[1245] = f[516] && !f[432] && !f[515] && f[380]; // c6t936i93
	assign leaf[1246] = f[516] && !f[432] && f[515] && !f[462]; // c6t936i93
	assign leaf[1247] = f[516] && !f[432] && f[515] && f[462]; // c6t936i93
	assign leaf[1248] = f[516] && f[432] && !f[155] && !f[209]; // c6t936i93
	assign leaf[1249] = f[516] && f[432] && !f[155] && f[209]; // c6t936i93
	assign leaf[1250] = f[516] && f[432] && f[155] && !f[573]; // c6t936i93
	assign leaf[1251] = f[516] && f[432] && f[155] && f[573]; // c6t936i93
	assign leaf[1252] = !f[656] && !f[146] && !f[351] && !f[299]; // c6t946i94
	assign leaf[1253] = !f[656] && !f[146] && !f[351] && f[299]; // c6t946i94
	assign leaf[1254] = !f[656] && !f[146] && f[351] && !f[491]; // c6t946i94
	assign leaf[1255] = !f[656] && !f[146] && f[351] && f[491]; // c6t946i94
	assign leaf[1256] = !f[656] && f[146]; // c6t946i94
	assign leaf[1257] = f[656] && !f[181] && !f[157] && !f[266]; // c6t946i94
	assign leaf[1258] = f[656] && !f[181] && !f[157] && f[266]; // c6t946i94
	assign leaf[1259] = f[656] && !f[181] && f[157] && !f[242]; // c6t946i94
	assign leaf[1260] = f[656] && !f[181] && f[157] && f[242]; // c6t946i94
	assign leaf[1261] = f[656] && f[181] && !f[605]; // c6t946i94
	assign leaf[1262] = f[656] && f[181] && f[605] && !f[578]; // c6t946i94
	assign leaf[1263] = f[656] && f[181] && f[605] && f[578]; // c6t946i94
	assign leaf[1264] = !f[661] && !f[262] && !f[521] && !f[490]; // c6t956i95
	assign leaf[1265] = !f[661] && !f[262] && !f[521] && f[490]; // c6t956i95
	assign leaf[1266] = !f[661] && !f[262] && f[521] && !f[348]; // c6t956i95
	assign leaf[1267] = !f[661] && !f[262] && f[521] && f[348]; // c6t956i95
	assign leaf[1268] = !f[661] && f[262] && !f[124] && !f[568]; // c6t956i95
	assign leaf[1269] = !f[661] && f[262] && !f[124] && f[568]; // c6t956i95
	assign leaf[1270] = !f[661] && f[262] && f[124] && !f[156]; // c6t956i95
	assign leaf[1271] = !f[661] && f[262] && f[124] && f[156]; // c6t956i95
	assign leaf[1272] = f[661] && !f[552] && !f[321] && !f[237]; // c6t956i95
	assign leaf[1273] = f[661] && !f[552] && !f[321] && f[237]; // c6t956i95
	assign leaf[1274] = f[661] && !f[552] && f[321]; // c6t956i95
	assign leaf[1275] = f[661] && f[552] && !f[233] && !f[234]; // c6t956i95
	assign leaf[1276] = f[661] && f[552] && !f[233] && f[234]; // c6t956i95
	assign leaf[1277] = f[661] && f[552] && f[233] && !f[128]; // c6t956i95
	assign leaf[1278] = f[661] && f[552] && f[233] && f[128]; // c6t956i95
	assign leaf[1279] = !f[267] && !f[120] && !f[237] && !f[155]; // c6t966i96
	assign leaf[1280] = !f[267] && !f[120] && !f[237] && f[155]; // c6t966i96
	assign leaf[1281] = !f[267] && !f[120] && f[237] && !f[634]; // c6t966i96
	assign leaf[1282] = !f[267] && !f[120] && f[237] && f[634]; // c6t966i96
	assign leaf[1283] = !f[267] && f[120]; // c6t966i96
	assign leaf[1284] = f[267] && !f[321] && !f[659] && !f[551]; // c6t966i96
	assign leaf[1285] = f[267] && !f[321] && !f[659] && f[551]; // c6t966i96
	assign leaf[1286] = f[267] && !f[321] && f[659]; // c6t966i96
	assign leaf[1287] = f[267] && f[321] && !f[181] && !f[433]; // c6t966i96
	assign leaf[1288] = f[267] && f[321] && !f[181] && f[433]; // c6t966i96
	assign leaf[1289] = f[267] && f[321] && f[181] && !f[495]; // c6t966i96
	assign leaf[1290] = f[267] && f[321] && f[181] && f[495]; // c6t966i96
	assign leaf[1291] = !f[547] && !f[631] && !f[603] && !f[463]; // c6t976i97
	assign leaf[1292] = !f[547] && !f[631] && !f[603] && f[463]; // c6t976i97
	assign leaf[1293] = !f[547] && !f[631] && f[603] && !f[493]; // c6t976i97
	assign leaf[1294] = !f[547] && !f[631] && f[603] && f[493]; // c6t976i97
	assign leaf[1295] = !f[547] && f[631] && !f[178] && !f[267]; // c6t976i97
	assign leaf[1296] = !f[547] && f[631] && !f[178] && f[267]; // c6t976i97
	assign leaf[1297] = !f[547] && f[631] && f[178] && !f[456]; // c6t976i97
	assign leaf[1298] = !f[547] && f[631] && f[178] && f[456]; // c6t976i97
	assign leaf[1299] = f[547] && !f[488] && !f[572] && !f[513]; // c6t976i97
	assign leaf[1300] = f[547] && !f[488] && !f[572] && f[513]; // c6t976i97
	assign leaf[1301] = f[547] && !f[488] && f[572] && !f[154]; // c6t976i97
	assign leaf[1302] = f[547] && !f[488] && f[572] && f[154]; // c6t976i97
	assign leaf[1303] = f[547] && f[488] && !f[631] && !f[514]; // c6t976i97
	assign leaf[1304] = f[547] && f[488] && !f[631] && f[514]; // c6t976i97
	assign leaf[1305] = f[547] && f[488] && f[631] && !f[573]; // c6t976i97
	assign leaf[1306] = f[547] && f[488] && f[631] && f[573]; // c6t976i97
	assign leaf[1307] = !f[516] && !f[405] && !f[240] && !f[123]; // c6t986i98
	assign leaf[1308] = !f[516] && !f[405] && !f[240] && f[123]; // c6t986i98
	assign leaf[1309] = !f[516] && !f[405] && f[240] && !f[433]; // c6t986i98
	assign leaf[1310] = !f[516] && !f[405] && f[240] && f[433]; // c6t986i98
	assign leaf[1311] = !f[516] && f[405] && !f[486] && !f[455]; // c6t986i98
	assign leaf[1312] = !f[516] && f[405] && !f[486] && f[455]; // c6t986i98
	assign leaf[1313] = !f[516] && f[405] && f[486] && !f[233]; // c6t986i98
	assign leaf[1314] = !f[516] && f[405] && f[486] && f[233]; // c6t986i98
	assign leaf[1315] = f[516] && !f[432] && !f[486] && !f[377]; // c6t986i98
	assign leaf[1316] = f[516] && !f[432] && !f[486] && f[377]; // c6t986i98
	assign leaf[1317] = f[516] && !f[432] && f[486] && !f[631]; // c6t986i98
	assign leaf[1318] = f[516] && !f[432] && f[486] && f[631]; // c6t986i98
	assign leaf[1319] = f[516] && f[432] && !f[434] && !f[633]; // c6t986i98
	assign leaf[1320] = f[516] && f[432] && !f[434] && f[633]; // c6t986i98
	assign leaf[1321] = f[516] && f[432] && f[434] && !f[216]; // c6t986i98
	assign leaf[1322] = f[516] && f[432] && f[434] && f[216]; // c6t986i98
	assign leaf[1323] = !f[516] && !f[544] && !f[570] && !f[568]; // c6t996i99
	assign leaf[1324] = !f[516] && !f[544] && !f[570] && f[568]; // c6t996i99
	assign leaf[1325] = !f[516] && !f[544] && f[570] && !f[654]; // c6t996i99
	assign leaf[1326] = !f[516] && !f[544] && f[570] && f[654]; // c6t996i99
	assign leaf[1327] = !f[516] && f[544] && !f[457] && !f[320]; // c6t996i99
	assign leaf[1328] = !f[516] && f[544] && !f[457] && f[320]; // c6t996i99
	assign leaf[1329] = !f[516] && f[544] && f[457] && !f[373]; // c6t996i99
	assign leaf[1330] = !f[516] && f[544] && f[457] && f[373]; // c6t996i99
	assign leaf[1331] = f[516] && !f[601] && !f[660] && !f[295]; // c6t996i99
	assign leaf[1332] = f[516] && !f[601] && !f[660] && f[295]; // c6t996i99
	assign leaf[1333] = f[516] && !f[601] && f[660]; // c6t996i99
	assign leaf[1334] = f[516] && f[601] && !f[544]; // c6t996i99
	assign leaf[1335] = f[516] && f[601] && f[544] && !f[492]; // c6t996i99
	assign leaf[1336] = f[516] && f[601] && f[544] && f[492]; // c6t996i99
endmodule

module decision_tree_leaves_7(input logic [0:783] f, output logic [0:1279] leaf);
	assign leaf[0] = !f[739] && !f[742] && !f[709] && !f[712]; // c7t7i0
	assign leaf[1] = !f[739] && !f[742] && !f[709] && f[712]; // c7t7i0
	assign leaf[2] = !f[739] && !f[742] && f[709] && !f[405]; // c7t7i0
	assign leaf[3] = !f[739] && !f[742] && f[709] && f[405]; // c7t7i0
	assign leaf[4] = !f[739] && f[742] && !f[431] && !f[404]; // c7t7i0
	assign leaf[5] = !f[739] && f[742] && !f[431] && f[404]; // c7t7i0
	assign leaf[6] = !f[739] && f[742] && f[431] && !f[231]; // c7t7i0
	assign leaf[7] = !f[739] && f[742] && f[431] && f[231]; // c7t7i0
	assign leaf[8] = f[739] && !f[405] && !f[460] && !f[377]; // c7t7i0
	assign leaf[9] = f[739] && !f[405] && !f[460] && f[377]; // c7t7i0
	assign leaf[10] = f[739] && !f[405] && f[460] && !f[232]; // c7t7i0
	assign leaf[11] = f[739] && !f[405] && f[460] && f[232]; // c7t7i0
	assign leaf[12] = f[739] && f[405] && !f[233] && !f[207]; // c7t7i0
	assign leaf[13] = f[739] && f[405] && !f[233] && f[207]; // c7t7i0
	assign leaf[14] = f[739] && f[405] && f[233] && !f[374]; // c7t7i0
	assign leaf[15] = f[739] && f[405] && f[233] && f[374]; // c7t7i0
	assign leaf[16] = !f[405] && !f[155] && !f[457] && !f[568]; // c7t17i1
	assign leaf[17] = !f[405] && !f[155] && !f[457] && f[568]; // c7t17i1
	assign leaf[18] = !f[405] && !f[155] && f[457] && !f[229]; // c7t17i1
	assign leaf[19] = !f[405] && !f[155] && f[457] && f[229]; // c7t17i1
	assign leaf[20] = !f[405] && f[155] && !f[678] && !f[578]; // c7t17i1
	assign leaf[21] = !f[405] && f[155] && !f[678] && f[578]; // c7t17i1
	assign leaf[22] = !f[405] && f[155] && f[678] && !f[603]; // c7t17i1
	assign leaf[23] = !f[405] && f[155] && f[678] && f[603]; // c7t17i1
	assign leaf[24] = f[405] && !f[231] && !f[708] && !f[710]; // c7t17i1
	assign leaf[25] = f[405] && !f[231] && !f[708] && f[710]; // c7t17i1
	assign leaf[26] = f[405] && !f[231] && f[708] && !f[542]; // c7t17i1
	assign leaf[27] = f[405] && !f[231] && f[708] && f[542]; // c7t17i1
	assign leaf[28] = f[405] && f[231] && !f[606] && !f[264]; // c7t17i1
	assign leaf[29] = f[405] && f[231] && !f[606] && f[264]; // c7t17i1
	assign leaf[30] = f[405] && f[231] && f[606] && !f[312]; // c7t17i1
	assign leaf[31] = f[405] && f[231] && f[606] && f[312]; // c7t17i1
	assign leaf[32] = !f[405] && !f[156] && !f[458] && !f[153]; // c7t27i2
	assign leaf[33] = !f[405] && !f[156] && !f[458] && f[153]; // c7t27i2
	assign leaf[34] = !f[405] && !f[156] && f[458] && !f[231]; // c7t27i2
	assign leaf[35] = !f[405] && !f[156] && f[458] && f[231]; // c7t27i2
	assign leaf[36] = !f[405] && f[156] && !f[678] && !f[597]; // c7t27i2
	assign leaf[37] = !f[405] && f[156] && !f[678] && f[597]; // c7t27i2
	assign leaf[38] = !f[405] && f[156] && f[678] && !f[570]; // c7t27i2
	assign leaf[39] = !f[405] && f[156] && f[678] && f[570]; // c7t27i2
	assign leaf[40] = f[405] && !f[231] && !f[257] && !f[705]; // c7t27i2
	assign leaf[41] = f[405] && !f[231] && !f[257] && f[705]; // c7t27i2
	assign leaf[42] = f[405] && !f[231] && f[257] && !f[289]; // c7t27i2
	assign leaf[43] = f[405] && !f[231] && f[257] && f[289]; // c7t27i2
	assign leaf[44] = f[405] && f[231] && !f[519] && !f[500]; // c7t27i2
	assign leaf[45] = f[405] && f[231] && !f[519] && f[500]; // c7t27i2
	assign leaf[46] = f[405] && f[231] && f[519] && !f[550]; // c7t27i2
	assign leaf[47] = f[405] && f[231] && f[519] && f[550]; // c7t27i2
	assign leaf[48] = !f[405] && !f[268] && !f[430] && !f[154]; // c7t37i3
	assign leaf[49] = !f[405] && !f[268] && !f[430] && f[154]; // c7t37i3
	assign leaf[50] = !f[405] && !f[268] && f[430] && !f[256]; // c7t37i3
	assign leaf[51] = !f[405] && !f[268] && f[430] && f[256]; // c7t37i3
	assign leaf[52] = !f[405] && f[268] && !f[156] && !f[430]; // c7t37i3
	assign leaf[53] = !f[405] && f[268] && !f[156] && f[430]; // c7t37i3
	assign leaf[54] = !f[405] && f[268] && f[156] && !f[490]; // c7t37i3
	assign leaf[55] = !f[405] && f[268] && f[156] && f[490]; // c7t37i3
	assign leaf[56] = f[405] && !f[268] && !f[707] && !f[312]; // c7t37i3
	assign leaf[57] = f[405] && !f[268] && !f[707] && f[312]; // c7t37i3
	assign leaf[58] = f[405] && !f[268] && f[707] && !f[515]; // c7t37i3
	assign leaf[59] = f[405] && !f[268] && f[707] && f[515]; // c7t37i3
	assign leaf[60] = f[405] && f[268] && !f[235] && !f[285]; // c7t37i3
	assign leaf[61] = f[405] && f[268] && !f[235] && f[285]; // c7t37i3
	assign leaf[62] = f[405] && f[268] && f[235] && !f[376]; // c7t37i3
	assign leaf[63] = f[405] && f[268] && f[235] && f[376]; // c7t37i3
	assign leaf[64] = !f[404] && !f[155] && !f[428] && !f[377]; // c7t47i4
	assign leaf[65] = !f[404] && !f[155] && !f[428] && f[377]; // c7t47i4
	assign leaf[66] = !f[404] && !f[155] && f[428] && !f[487]; // c7t47i4
	assign leaf[67] = !f[404] && !f[155] && f[428] && f[487]; // c7t47i4
	assign leaf[68] = !f[404] && f[155] && !f[678] && !f[127]; // c7t47i4
	assign leaf[69] = !f[404] && f[155] && !f[678] && f[127]; // c7t47i4
	assign leaf[70] = !f[404] && f[155] && f[678] && !f[603]; // c7t47i4
	assign leaf[71] = !f[404] && f[155] && f[678] && f[603]; // c7t47i4
	assign leaf[72] = f[404] && !f[412] && !f[441] && !f[345]; // c7t47i4
	assign leaf[73] = f[404] && !f[412] && !f[441] && f[345]; // c7t47i4
	assign leaf[74] = f[404] && !f[412] && f[441] && !f[714]; // c7t47i4
	assign leaf[75] = f[404] && !f[412] && f[441] && f[714]; // c7t47i4
	assign leaf[76] = f[404] && f[412] && !f[715] && !f[710]; // c7t47i4
	assign leaf[77] = f[404] && f[412] && !f[715] && f[710]; // c7t47i4
	assign leaf[78] = f[404] && f[412] && f[715] && !f[322]; // c7t47i4
	assign leaf[79] = f[404] && f[412] && f[715] && f[322]; // c7t47i4
	assign leaf[80] = !f[404] && !f[157] && !f[269] && !f[461]; // c7t57i5
	assign leaf[81] = !f[404] && !f[157] && !f[269] && f[461]; // c7t57i5
	assign leaf[82] = !f[404] && !f[157] && f[269] && !f[541]; // c7t57i5
	assign leaf[83] = !f[404] && !f[157] && f[269] && f[541]; // c7t57i5
	assign leaf[84] = !f[404] && f[157] && !f[203] && !f[679]; // c7t57i5
	assign leaf[85] = !f[404] && f[157] && !f[203] && f[679]; // c7t57i5
	assign leaf[86] = !f[404] && f[157] && f[203] && !f[606]; // c7t57i5
	assign leaf[87] = !f[404] && f[157] && f[203] && f[606]; // c7t57i5
	assign leaf[88] = f[404] && !f[155] && !f[412] && !f[296]; // c7t57i5
	assign leaf[89] = f[404] && !f[155] && !f[412] && f[296]; // c7t57i5
	assign leaf[90] = f[404] && !f[155] && f[412] && !f[323]; // c7t57i5
	assign leaf[91] = f[404] && !f[155] && f[412] && f[323]; // c7t57i5
	assign leaf[92] = f[404] && f[155]; // c7t57i5
	assign leaf[93] = !f[377] && !f[459] && !f[512] && !f[158]; // c7t67i6
	assign leaf[94] = !f[377] && !f[459] && !f[512] && f[158]; // c7t67i6
	assign leaf[95] = !f[377] && !f[459] && f[512] && !f[715]; // c7t67i6
	assign leaf[96] = !f[377] && !f[459] && f[512] && f[715]; // c7t67i6
	assign leaf[97] = !f[377] && f[459] && !f[373] && !f[324]; // c7t67i6
	assign leaf[98] = !f[377] && f[459] && !f[373] && f[324]; // c7t67i6
	assign leaf[99] = !f[377] && f[459] && f[373] && !f[285]; // c7t67i6
	assign leaf[100] = !f[377] && f[459] && f[373] && f[285]; // c7t67i6
	assign leaf[101] = f[377] && !f[339] && !f[385] && !f[517]; // c7t67i6
	assign leaf[102] = f[377] && !f[339] && !f[385] && f[517]; // c7t67i6
	assign leaf[103] = f[377] && !f[339] && f[385] && !f[186]; // c7t67i6
	assign leaf[104] = f[377] && !f[339] && f[385] && f[186]; // c7t67i6
	assign leaf[105] = f[377] && f[339] && !f[257] && !f[269]; // c7t67i6
	assign leaf[106] = f[377] && f[339] && !f[257] && f[269]; // c7t67i6
	assign leaf[107] = f[377] && f[339] && f[257]; // c7t67i6
	assign leaf[108] = !f[154] && !f[432] && !f[513] && !f[378]; // c7t77i7
	assign leaf[109] = !f[154] && !f[432] && !f[513] && f[378]; // c7t77i7
	assign leaf[110] = !f[154] && !f[432] && f[513] && !f[399]; // c7t77i7
	assign leaf[111] = !f[154] && !f[432] && f[513] && f[399]; // c7t77i7
	assign leaf[112] = !f[154] && f[432] && !f[232] && !f[205]; // c7t77i7
	assign leaf[113] = !f[154] && f[432] && !f[232] && f[205]; // c7t77i7
	assign leaf[114] = !f[154] && f[432] && f[232] && !f[578]; // c7t77i7
	assign leaf[115] = !f[154] && f[432] && f[232] && f[578]; // c7t77i7
	assign leaf[116] = f[154] && !f[577] && !f[679] && !f[296]; // c7t77i7
	assign leaf[117] = f[154] && !f[577] && !f[679] && f[296]; // c7t77i7
	assign leaf[118] = f[154] && !f[577] && f[679] && !f[571]; // c7t77i7
	assign leaf[119] = f[154] && !f[577] && f[679] && f[571]; // c7t77i7
	assign leaf[120] = f[154] && f[577] && !f[284] && !f[145]; // c7t77i7
	assign leaf[121] = f[154] && f[577] && !f[284] && f[145]; // c7t77i7
	assign leaf[122] = f[154] && f[577] && f[284]; // c7t77i7
	assign leaf[123] = !f[267] && !f[745] && !f[402] && !f[377]; // c7t87i8
	assign leaf[124] = !f[267] && !f[745] && !f[402] && f[377]; // c7t87i8
	assign leaf[125] = !f[267] && !f[745] && f[402] && !f[295]; // c7t87i8
	assign leaf[126] = !f[267] && !f[745] && f[402] && f[295]; // c7t87i8
	assign leaf[127] = !f[267] && f[745] && !f[432] && !f[373]; // c7t87i8
	assign leaf[128] = !f[267] && f[745] && !f[432] && f[373]; // c7t87i8
	assign leaf[129] = !f[267] && f[745] && f[432]; // c7t87i8
	assign leaf[130] = f[267] && !f[263] && !f[236] && !f[290]; // c7t87i8
	assign leaf[131] = f[267] && !f[263] && !f[236] && f[290]; // c7t87i8
	assign leaf[132] = f[267] && !f[263] && f[236] && !f[606]; // c7t87i8
	assign leaf[133] = f[267] && !f[263] && f[236] && f[606]; // c7t87i8
	assign leaf[134] = f[267] && f[263] && !f[567] && !f[403]; // c7t87i8
	assign leaf[135] = f[267] && f[263] && !f[567] && f[403]; // c7t87i8
	assign leaf[136] = f[267] && f[263] && f[567] && !f[677]; // c7t87i8
	assign leaf[137] = f[267] && f[263] && f[567] && f[677]; // c7t87i8
	assign leaf[138] = !f[157] && !f[376] && !f[552] && !f[401]; // c7t97i9
	assign leaf[139] = !f[157] && !f[376] && !f[552] && f[401]; // c7t97i9
	assign leaf[140] = !f[157] && !f[376] && f[552] && !f[746]; // c7t97i9
	assign leaf[141] = !f[157] && !f[376] && f[552] && f[746]; // c7t97i9
	assign leaf[142] = !f[157] && f[376] && !f[340] && !f[411]; // c7t97i9
	assign leaf[143] = !f[157] && f[376] && !f[340] && f[411]; // c7t97i9
	assign leaf[144] = !f[157] && f[376] && f[340] && !f[430]; // c7t97i9
	assign leaf[145] = !f[157] && f[376] && f[340] && f[430]; // c7t97i9
	assign leaf[146] = f[157] && !f[518]; // c7t97i9
	assign leaf[147] = f[157] && f[518] && !f[148] && !f[685]; // c7t97i9
	assign leaf[148] = f[157] && f[518] && !f[148] && f[685]; // c7t97i9
	assign leaf[149] = f[157] && f[518] && f[148] && !f[552]; // c7t97i9
	assign leaf[150] = f[157] && f[518] && f[148] && f[552]; // c7t97i9
	assign leaf[151] = !f[154] && !f[159] && !f[432] && !f[486]; // c7t107i10
	assign leaf[152] = !f[154] && !f[159] && !f[432] && f[486]; // c7t107i10
	assign leaf[153] = !f[154] && !f[159] && f[432] && !f[345]; // c7t107i10
	assign leaf[154] = !f[154] && !f[159] && f[432] && f[345]; // c7t107i10
	assign leaf[155] = !f[154] && f[159] && !f[206]; // c7t107i10
	assign leaf[156] = !f[154] && f[159] && f[206] && !f[268]; // c7t107i10
	assign leaf[157] = !f[154] && f[159] && f[206] && f[268]; // c7t107i10
	assign leaf[158] = f[154] && !f[577] && !f[679] && !f[240]; // c7t107i10
	assign leaf[159] = f[154] && !f[577] && !f[679] && f[240]; // c7t107i10
	assign leaf[160] = f[154] && !f[577] && f[679] && !f[377]; // c7t107i10
	assign leaf[161] = f[154] && !f[577] && f[679] && f[377]; // c7t107i10
	assign leaf[162] = f[154] && f[577] && !f[145]; // c7t107i10
	assign leaf[163] = f[154] && f[577] && f[145]; // c7t107i10
	assign leaf[164] = !f[376] && !f[297] && !f[707] && !f[232]; // c7t117i11
	assign leaf[165] = !f[376] && !f[297] && !f[707] && f[232]; // c7t117i11
	assign leaf[166] = !f[376] && !f[297] && f[707] && !f[243]; // c7t117i11
	assign leaf[167] = !f[376] && !f[297] && f[707] && f[243]; // c7t117i11
	assign leaf[168] = !f[376] && f[297] && !f[266] && !f[607]; // c7t117i11
	assign leaf[169] = !f[376] && f[297] && !f[266] && f[607]; // c7t117i11
	assign leaf[170] = !f[376] && f[297] && f[266] && !f[581]; // c7t117i11
	assign leaf[171] = !f[376] && f[297] && f[266] && f[581]; // c7t117i11
	assign leaf[172] = f[376] && !f[312] && !f[184] && !f[355]; // c7t117i11
	assign leaf[173] = f[376] && !f[312] && !f[184] && f[355]; // c7t117i11
	assign leaf[174] = f[376] && !f[312] && f[184] && !f[347]; // c7t117i11
	assign leaf[175] = f[376] && !f[312] && f[184] && f[347]; // c7t117i11
	assign leaf[176] = f[376] && f[312] && !f[581] && !f[346]; // c7t117i11
	assign leaf[177] = f[376] && f[312] && !f[581] && f[346]; // c7t117i11
	assign leaf[178] = f[376] && f[312] && f[581] && !f[413]; // c7t117i11
	assign leaf[179] = f[376] && f[312] && f[581] && f[413]; // c7t117i11
	assign leaf[180] = !f[158] && !f[153] && !f[432] && !f[377]; // c7t127i12
	assign leaf[181] = !f[158] && !f[153] && !f[432] && f[377]; // c7t127i12
	assign leaf[182] = !f[158] && !f[153] && f[432] && !f[372]; // c7t127i12
	assign leaf[183] = !f[158] && !f[153] && f[432] && f[372]; // c7t127i12
	assign leaf[184] = !f[158] && f[153] && !f[604] && !f[634]; // c7t127i12
	assign leaf[185] = !f[158] && f[153] && !f[604] && f[634]; // c7t127i12
	assign leaf[186] = !f[158] && f[153] && f[604] && !f[687]; // c7t127i12
	assign leaf[187] = !f[158] && f[153] && f[604] && f[687]; // c7t127i12
	assign leaf[188] = f[158] && !f[686] && !f[149] && !f[687]; // c7t127i12
	assign leaf[189] = f[158] && !f[686] && !f[149] && f[687]; // c7t127i12
	assign leaf[190] = f[158] && !f[686] && f[149] && !f[605]; // c7t127i12
	assign leaf[191] = f[158] && !f[686] && f[149] && f[605]; // c7t127i12
	assign leaf[192] = f[158] && f[686] && !f[573]; // c7t127i12
	assign leaf[193] = f[158] && f[686] && f[573] && !f[374]; // c7t127i12
	assign leaf[194] = f[158] && f[686] && f[573] && f[374]; // c7t127i12
	assign leaf[195] = !f[569] && !f[267] && !f[433] && !f[487]; // c7t137i13
	assign leaf[196] = !f[569] && !f[267] && !f[433] && f[487]; // c7t137i13
	assign leaf[197] = !f[569] && !f[267] && f[433] && !f[346]; // c7t137i13
	assign leaf[198] = !f[569] && !f[267] && f[433] && f[346]; // c7t137i13
	assign leaf[199] = !f[569] && f[267] && !f[263] && !f[236]; // c7t137i13
	assign leaf[200] = !f[569] && f[267] && !f[263] && f[236]; // c7t137i13
	assign leaf[201] = !f[569] && f[267] && f[263] && !f[260]; // c7t137i13
	assign leaf[202] = !f[569] && f[267] && f[263] && f[260]; // c7t137i13
	assign leaf[203] = f[569] && !f[679] && !f[677] && !f[709]; // c7t137i13
	assign leaf[204] = f[569] && !f[679] && !f[677] && f[709]; // c7t137i13
	assign leaf[205] = f[569] && !f[679] && f[677] && !f[238]; // c7t137i13
	assign leaf[206] = f[569] && !f[679] && f[677] && f[238]; // c7t137i13
	assign leaf[207] = f[569] && f[679] && !f[271] && !f[326]; // c7t137i13
	assign leaf[208] = f[569] && f[679] && !f[271] && f[326]; // c7t137i13
	assign leaf[209] = f[569] && f[679] && f[271] && !f[602]; // c7t137i13
	assign leaf[210] = f[569] && f[679] && f[271] && f[602]; // c7t137i13
	assign leaf[211] = !f[580] && !f[259] && !f[206] && !f[459]; // c7t147i14
	assign leaf[212] = !f[580] && !f[259] && !f[206] && f[459]; // c7t147i14
	assign leaf[213] = !f[580] && !f[259] && f[206] && !f[578]; // c7t147i14
	assign leaf[214] = !f[580] && !f[259] && f[206] && f[578]; // c7t147i14
	assign leaf[215] = !f[580] && f[259] && !f[263] && !f[427]; // c7t147i14
	assign leaf[216] = !f[580] && f[259] && !f[263] && f[427]; // c7t147i14
	assign leaf[217] = !f[580] && f[259] && f[263] && !f[554]; // c7t147i14
	assign leaf[218] = !f[580] && f[259] && f[263] && f[554]; // c7t147i14
	assign leaf[219] = f[580] && !f[746] && !f[283] && !f[749]; // c7t147i14
	assign leaf[220] = f[580] && !f[746] && !f[283] && f[749]; // c7t147i14
	assign leaf[221] = f[580] && !f[746] && f[283] && !f[206]; // c7t147i14
	assign leaf[222] = f[580] && !f[746] && f[283] && f[206]; // c7t147i14
	assign leaf[223] = f[580] && f[746] && !f[436]; // c7t147i14
	assign leaf[224] = f[580] && f[746] && f[436]; // c7t147i14
	assign leaf[225] = !f[744] && !f[578] && !f[437] && !f[711]; // c7t157i15
	assign leaf[226] = !f[744] && !f[578] && !f[437] && f[711]; // c7t157i15
	assign leaf[227] = !f[744] && !f[578] && f[437] && !f[296]; // c7t157i15
	assign leaf[228] = !f[744] && !f[578] && f[437] && f[296]; // c7t157i15
	assign leaf[229] = !f[744] && f[578] && !f[717] && !f[340]; // c7t157i15
	assign leaf[230] = !f[744] && f[578] && !f[717] && f[340]; // c7t157i15
	assign leaf[231] = !f[744] && f[578] && f[717] && !f[460]; // c7t157i15
	assign leaf[232] = !f[744] && f[578] && f[717] && f[460]; // c7t157i15
	assign leaf[233] = f[744] && !f[461] && !f[349] && !f[374]; // c7t157i15
	assign leaf[234] = f[744] && !f[461] && !f[349] && f[374]; // c7t157i15
	assign leaf[235] = f[744] && !f[461] && f[349] && !f[238]; // c7t157i15
	assign leaf[236] = f[744] && !f[461] && f[349] && f[238]; // c7t157i15
	assign leaf[237] = f[744] && f[461] && !f[458] && !f[518]; // c7t157i15
	assign leaf[238] = f[744] && f[461] && !f[458] && f[518]; // c7t157i15
	assign leaf[239] = f[744] && f[461] && f[458] && !f[344]; // c7t157i15
	assign leaf[240] = f[744] && f[461] && f[458] && f[344]; // c7t157i15
	assign leaf[241] = !f[376] && !f[607] && !f[402] && !f[427]; // c7t167i16
	assign leaf[242] = !f[376] && !f[607] && !f[402] && f[427]; // c7t167i16
	assign leaf[243] = !f[376] && !f[607] && f[402] && !f[431]; // c7t167i16
	assign leaf[244] = !f[376] && !f[607] && f[402] && f[431]; // c7t167i16
	assign leaf[245] = !f[376] && f[607] && !f[435] && !f[717]; // c7t167i16
	assign leaf[246] = !f[376] && f[607] && !f[435] && f[717]; // c7t167i16
	assign leaf[247] = !f[376] && f[607] && f[435] && !f[227]; // c7t167i16
	assign leaf[248] = !f[376] && f[607] && f[435] && f[227]; // c7t167i16
	assign leaf[249] = f[376] && !f[384] && !f[410] && !f[740]; // c7t167i16
	assign leaf[250] = f[376] && !f[384] && !f[410] && f[740]; // c7t167i16
	assign leaf[251] = f[376] && !f[384] && f[410] && !f[349]; // c7t167i16
	assign leaf[252] = f[376] && !f[384] && f[410] && f[349]; // c7t167i16
	assign leaf[253] = f[376] && f[384] && !f[183] && !f[569]; // c7t167i16
	assign leaf[254] = f[376] && f[384] && !f[183] && f[569]; // c7t167i16
	assign leaf[255] = f[376] && f[384] && f[183] && !f[715]; // c7t167i16
	assign leaf[256] = f[376] && f[384] && f[183] && f[715]; // c7t167i16
	assign leaf[257] = !f[159] && !f[298] && !f[348] && !f[296]; // c7t177i17
	assign leaf[258] = !f[159] && !f[298] && !f[348] && f[296]; // c7t177i17
	assign leaf[259] = !f[159] && !f[298] && f[348] && !f[340]; // c7t177i17
	assign leaf[260] = !f[159] && !f[298] && f[348] && f[340]; // c7t177i17
	assign leaf[261] = !f[159] && f[298] && !f[266] && !f[294]; // c7t177i17
	assign leaf[262] = !f[159] && f[298] && !f[266] && f[294]; // c7t177i17
	assign leaf[263] = !f[159] && f[298] && f[266] && !f[553]; // c7t177i17
	assign leaf[264] = !f[159] && f[298] && f[266] && f[553]; // c7t177i17
	assign leaf[265] = f[159] && !f[149]; // c7t177i17
	assign leaf[266] = f[159] && f[149]; // c7t177i17
	assign leaf[267] = !f[348] && !f[239] && !f[321] && !f[486]; // c7t187i18
	assign leaf[268] = !f[348] && !f[239] && !f[321] && f[486]; // c7t187i18
	assign leaf[269] = !f[348] && !f[239] && f[321] && !f[182]; // c7t187i18
	assign leaf[270] = !f[348] && !f[239] && f[321] && f[182]; // c7t187i18
	assign leaf[271] = !f[348] && f[239] && !f[579] && !f[234]; // c7t187i18
	assign leaf[272] = !f[348] && f[239] && !f[579] && f[234]; // c7t187i18
	assign leaf[273] = !f[348] && f[239] && f[579] && !f[717]; // c7t187i18
	assign leaf[274] = !f[348] && f[239] && f[579] && f[717]; // c7t187i18
	assign leaf[275] = f[348] && !f[328] && !f[285] && !f[266]; // c7t187i18
	assign leaf[276] = f[348] && !f[328] && !f[285] && f[266]; // c7t187i18
	assign leaf[277] = f[348] && !f[328] && f[285] && !f[318]; // c7t187i18
	assign leaf[278] = f[348] && !f[328] && f[285] && f[318]; // c7t187i18
	assign leaf[279] = f[348] && f[328] && !f[184] && !f[432]; // c7t187i18
	assign leaf[280] = f[348] && f[328] && !f[184] && f[432]; // c7t187i18
	assign leaf[281] = f[348] && f[328] && f[184] && !f[350]; // c7t187i18
	assign leaf[282] = f[348] && f[328] && f[184] && f[350]; // c7t187i18
	assign leaf[283] = !f[539] && !f[608] && !f[267] && !f[434]; // c7t197i19
	assign leaf[284] = !f[539] && !f[608] && !f[267] && f[434]; // c7t197i19
	assign leaf[285] = !f[539] && !f[608] && f[267] && !f[264]; // c7t197i19
	assign leaf[286] = !f[539] && !f[608] && f[267] && f[264]; // c7t197i19
	assign leaf[287] = !f[539] && f[608] && !f[746] && !f[210]; // c7t197i19
	assign leaf[288] = !f[539] && f[608] && !f[746] && f[210]; // c7t197i19
	assign leaf[289] = !f[539] && f[608] && f[746] && !f[207]; // c7t197i19
	assign leaf[290] = !f[539] && f[608] && f[746] && f[207]; // c7t197i19
	assign leaf[291] = f[539] && !f[714] && !f[229] && !f[712]; // c7t197i19
	assign leaf[292] = f[539] && !f[714] && !f[229] && f[712]; // c7t197i19
	assign leaf[293] = f[539] && !f[714] && f[229] && !f[569]; // c7t197i19
	assign leaf[294] = f[539] && !f[714] && f[229] && f[569]; // c7t197i19
	assign leaf[295] = f[539] && f[714] && !f[318]; // c7t197i19
	assign leaf[296] = f[539] && f[714] && f[318]; // c7t197i19
	assign leaf[297] = !f[376] && !f[461] && !f[515] && !f[406]; // c7t207i20
	assign leaf[298] = !f[376] && !f[461] && !f[515] && f[406]; // c7t207i20
	assign leaf[299] = !f[376] && !f[461] && f[515] && !f[484]; // c7t207i20
	assign leaf[300] = !f[376] && !f[461] && f[515] && f[484]; // c7t207i20
	assign leaf[301] = !f[376] && f[461] && !f[372] && !f[374]; // c7t207i20
	assign leaf[302] = !f[376] && f[461] && !f[372] && f[374]; // c7t207i20
	assign leaf[303] = !f[376] && f[461] && f[372] && !f[708]; // c7t207i20
	assign leaf[304] = !f[376] && f[461] && f[372] && f[708]; // c7t207i20
	assign leaf[305] = f[376] && !f[284] && !f[295] && !f[397]; // c7t207i20
	assign leaf[306] = f[376] && !f[284] && !f[295] && f[397]; // c7t207i20
	assign leaf[307] = f[376] && !f[284] && f[295] && !f[383]; // c7t207i20
	assign leaf[308] = f[376] && !f[284] && f[295] && f[383]; // c7t207i20
	assign leaf[309] = f[376] && f[284] && !f[553] && !f[271]; // c7t207i20
	assign leaf[310] = f[376] && f[284] && !f[553] && f[271]; // c7t207i20
	assign leaf[311] = f[376] && f[284] && f[553]; // c7t207i20
	assign leaf[312] = !f[566] && !f[270] && !f[324] && !f[678]; // c7t217i21
	assign leaf[313] = !f[566] && !f[270] && !f[324] && f[678]; // c7t217i21
	assign leaf[314] = !f[566] && !f[270] && f[324] && !f[570]; // c7t217i21
	assign leaf[315] = !f[566] && !f[270] && f[324] && f[570]; // c7t217i21
	assign leaf[316] = !f[566] && f[270] && !f[486] && !f[378]; // c7t217i21
	assign leaf[317] = !f[566] && f[270] && !f[486] && f[378]; // c7t217i21
	assign leaf[318] = !f[566] && f[270] && f[486] && !f[399]; // c7t217i21
	assign leaf[319] = !f[566] && f[270] && f[486] && f[399]; // c7t217i21
	assign leaf[320] = f[566] && !f[648] && !f[341] && !f[123]; // c7t217i21
	assign leaf[321] = f[566] && !f[648] && !f[341] && f[123]; // c7t217i21
	assign leaf[322] = f[566] && !f[648] && f[341]; // c7t217i21
	assign leaf[323] = f[566] && f[648]; // c7t217i21
	assign leaf[324] = !f[437] && !f[431] && !f[744] && !f[707]; // c7t227i22
	assign leaf[325] = !f[437] && !f[431] && !f[744] && f[707]; // c7t227i22
	assign leaf[326] = !f[437] && !f[431] && f[744] && !f[350]; // c7t227i22
	assign leaf[327] = !f[437] && !f[431] && f[744] && f[350]; // c7t227i22
	assign leaf[328] = !f[437] && f[431] && !f[466] && !f[383]; // c7t227i22
	assign leaf[329] = !f[437] && f[431] && !f[466] && f[383]; // c7t227i22
	assign leaf[330] = !f[437] && f[431] && f[466] && !f[411]; // c7t227i22
	assign leaf[331] = !f[437] && f[431] && f[466] && f[411]; // c7t227i22
	assign leaf[332] = f[437] && !f[606] && !f[232] && !f[484]; // c7t227i22
	assign leaf[333] = f[437] && !f[606] && !f[232] && f[484]; // c7t227i22
	assign leaf[334] = f[437] && !f[606] && f[232] && !f[343]; // c7t227i22
	assign leaf[335] = f[437] && !f[606] && f[232] && f[343]; // c7t227i22
	assign leaf[336] = f[437] && f[606] && !f[717] && !f[284]; // c7t227i22
	assign leaf[337] = f[437] && f[606] && !f[717] && f[284]; // c7t227i22
	assign leaf[338] = f[437] && f[606] && f[717] && !f[516]; // c7t227i22
	assign leaf[339] = f[437] && f[606] && f[717] && f[516]; // c7t227i22
	assign leaf[340] = !f[554] && !f[160] && !f[127] && !f[285]; // c7t237i23
	assign leaf[341] = !f[554] && !f[160] && !f[127] && f[285]; // c7t237i23
	assign leaf[342] = !f[554] && !f[160] && f[127] && !f[553]; // c7t237i23
	assign leaf[343] = !f[554] && !f[160] && f[127] && f[553]; // c7t237i23
	assign leaf[344] = !f[554] && f[160] && !f[152]; // c7t237i23
	assign leaf[345] = !f[554] && f[160] && f[152]; // c7t237i23
	assign leaf[346] = f[554] && !f[274] && !f[146] && !f[216]; // c7t237i23
	assign leaf[347] = f[554] && !f[274] && !f[146] && f[216]; // c7t237i23
	assign leaf[348] = f[554] && !f[274] && f[146]; // c7t237i23
	assign leaf[349] = f[554] && f[274]; // c7t237i23
	assign leaf[350] = !f[298] && !f[347] && !f[687] && !f[685]; // c7t247i24
	assign leaf[351] = !f[298] && !f[347] && !f[687] && f[685]; // c7t247i24
	assign leaf[352] = !f[298] && !f[347] && f[687] && !f[574]; // c7t247i24
	assign leaf[353] = !f[298] && !f[347] && f[687] && f[574]; // c7t247i24
	assign leaf[354] = !f[298] && f[347] && !f[341] && !f[355]; // c7t247i24
	assign leaf[355] = !f[298] && f[347] && !f[341] && f[355]; // c7t247i24
	assign leaf[356] = !f[298] && f[347] && f[341] && !f[240]; // c7t247i24
	assign leaf[357] = !f[298] && f[347] && f[341] && f[240]; // c7t247i24
	assign leaf[358] = f[298] && !f[182] && !f[460] && !f[542]; // c7t247i24
	assign leaf[359] = f[298] && !f[182] && !f[460] && f[542]; // c7t247i24
	assign leaf[360] = f[298] && !f[182] && f[460] && !f[400]; // c7t247i24
	assign leaf[361] = f[298] && !f[182] && f[460] && f[400]; // c7t247i24
	assign leaf[362] = f[298] && f[182] && !f[633] && !f[576]; // c7t247i24
	assign leaf[363] = f[298] && f[182] && !f[633] && f[576]; // c7t247i24
	assign leaf[364] = f[298] && f[182] && f[633] && !f[716]; // c7t247i24
	assign leaf[365] = f[298] && f[182] && f[633] && f[716]; // c7t247i24
	assign leaf[366] = !f[607] && !f[438] && !f[349] && !f[432]; // c7t257i25
	assign leaf[367] = !f[607] && !f[438] && !f[349] && f[432]; // c7t257i25
	assign leaf[368] = !f[607] && !f[438] && f[349] && !f[294]; // c7t257i25
	assign leaf[369] = !f[607] && !f[438] && f[349] && f[294]; // c7t257i25
	assign leaf[370] = !f[607] && f[438] && !f[540] && !f[372]; // c7t257i25
	assign leaf[371] = !f[607] && f[438] && !f[540] && f[372]; // c7t257i25
	assign leaf[372] = !f[607] && f[438] && f[540] && !f[233]; // c7t257i25
	assign leaf[373] = !f[607] && f[438] && f[540] && f[233]; // c7t257i25
	assign leaf[374] = f[607] && !f[435] && !f[180] && !f[319]; // c7t257i25
	assign leaf[375] = f[607] && !f[435] && !f[180] && f[319]; // c7t257i25
	assign leaf[376] = f[607] && !f[435] && f[180] && !f[173]; // c7t257i25
	assign leaf[377] = f[607] && !f[435] && f[180] && f[173]; // c7t257i25
	assign leaf[378] = f[607] && f[435] && !f[228] && !f[718]; // c7t257i25
	assign leaf[379] = f[607] && f[435] && !f[228] && f[718]; // c7t257i25
	assign leaf[380] = f[607] && f[435] && f[228] && !f[261]; // c7t257i25
	assign leaf[381] = f[607] && f[435] && f[228] && f[261]; // c7t257i25
	assign leaf[382] = !f[159] && !f[124] && !f[582] && !f[349]; // c7t267i26
	assign leaf[383] = !f[159] && !f[124] && !f[582] && f[349]; // c7t267i26
	assign leaf[384] = !f[159] && !f[124] && f[582] && !f[722]; // c7t267i26
	assign leaf[385] = !f[159] && !f[124] && f[582] && f[722]; // c7t267i26
	assign leaf[386] = !f[159] && f[124] && !f[399]; // c7t267i26
	assign leaf[387] = !f[159] && f[124] && f[399]; // c7t267i26
	assign leaf[388] = f[159] && !f[205] && !f[679]; // c7t267i26
	assign leaf[389] = f[159] && !f[205] && f[679] && !f[487]; // c7t267i26
	assign leaf[390] = f[159] && !f[205] && f[679] && f[487]; // c7t267i26
	assign leaf[391] = f[159] && f[205] && !f[297]; // c7t267i26
	assign leaf[392] = f[159] && f[205] && f[297]; // c7t267i26
	assign leaf[393] = !f[581] && !f[566] && !f[128] && !f[240]; // c7t277i27
	assign leaf[394] = !f[581] && !f[566] && !f[128] && f[240]; // c7t277i27
	assign leaf[395] = !f[581] && !f[566] && f[128]; // c7t277i27
	assign leaf[396] = !f[581] && f[566] && !f[620] && !f[178]; // c7t277i27
	assign leaf[397] = !f[581] && f[566] && !f[620] && f[178]; // c7t277i27
	assign leaf[398] = !f[581] && f[566] && f[620]; // c7t277i27
	assign leaf[399] = f[581] && !f[292] && !f[127] && !f[721]; // c7t277i27
	assign leaf[400] = f[581] && !f[292] && !f[127] && f[721]; // c7t277i27
	assign leaf[401] = f[581] && !f[292] && f[127]; // c7t277i27
	assign leaf[402] = f[581] && f[292] && !f[603] && !f[437]; // c7t277i27
	assign leaf[403] = f[581] && f[292] && !f[603] && f[437]; // c7t277i27
	assign leaf[404] = f[581] && f[292] && f[603] && !f[573]; // c7t277i27
	assign leaf[405] = f[581] && f[292] && f[603] && f[573]; // c7t277i27
	assign leaf[406] = !f[124] && !f[161] && !f[527] && !f[266]; // c7t287i28
	assign leaf[407] = !f[124] && !f[161] && !f[527] && f[266]; // c7t287i28
	assign leaf[408] = !f[124] && !f[161] && f[527] && !f[511]; // c7t287i28
	assign leaf[409] = !f[124] && !f[161] && f[527] && f[511]; // c7t287i28
	assign leaf[410] = !f[124] && f[161] && !f[178]; // c7t287i28
	assign leaf[411] = !f[124] && f[161] && f[178]; // c7t287i28
	assign leaf[412] = f[124] && !f[427]; // c7t287i28
	assign leaf[413] = f[124] && f[427]; // c7t287i28
	assign leaf[414] = !f[744] && !f[577] && !f[662] && !f[207]; // c7t297i29
	assign leaf[415] = !f[744] && !f[577] && !f[662] && f[207]; // c7t297i29
	assign leaf[416] = !f[744] && !f[577] && f[662] && !f[178]; // c7t297i29
	assign leaf[417] = !f[744] && !f[577] && f[662] && f[178]; // c7t297i29
	assign leaf[418] = !f[744] && f[577] && !f[655] && !f[489]; // c7t297i29
	assign leaf[419] = !f[744] && f[577] && !f[655] && f[489]; // c7t297i29
	assign leaf[420] = !f[744] && f[577] && f[655] && !f[573]; // c7t297i29
	assign leaf[421] = !f[744] && f[577] && f[655] && f[573]; // c7t297i29
	assign leaf[422] = f[744] && !f[433] && !f[488] && !f[349]; // c7t297i29
	assign leaf[423] = f[744] && !f[433] && !f[488] && f[349]; // c7t297i29
	assign leaf[424] = f[744] && !f[433] && f[488] && !f[260]; // c7t297i29
	assign leaf[425] = f[744] && !f[433] && f[488] && f[260]; // c7t297i29
	assign leaf[426] = f[744] && f[433] && !f[440] && !f[294]; // c7t297i29
	assign leaf[427] = f[744] && f[433] && !f[440] && f[294]; // c7t297i29
	assign leaf[428] = f[744] && f[433] && f[440]; // c7t297i29
	assign leaf[429] = !f[160] && !f[326] && !f[347] && !f[379]; // c7t307i30
	assign leaf[430] = !f[160] && !f[326] && !f[347] && f[379]; // c7t307i30
	assign leaf[431] = !f[160] && !f[326] && f[347] && !f[300]; // c7t307i30
	assign leaf[432] = !f[160] && !f[326] && f[347] && f[300]; // c7t307i30
	assign leaf[433] = !f[160] && f[326] && !f[433] && !f[488]; // c7t307i30
	assign leaf[434] = !f[160] && f[326] && !f[433] && f[488]; // c7t307i30
	assign leaf[435] = !f[160] && f[326] && f[433] && !f[489]; // c7t307i30
	assign leaf[436] = !f[160] && f[326] && f[433] && f[489]; // c7t307i30
	assign leaf[437] = f[160] && !f[687]; // c7t307i30
	assign leaf[438] = f[160] && f[687]; // c7t307i30
	assign leaf[439] = !f[677] && !f[595] && !f[542] && !f[294]; // c7t317i31
	assign leaf[440] = !f[677] && !f[595] && !f[542] && f[294]; // c7t317i31
	assign leaf[441] = !f[677] && !f[595] && f[542] && !f[241]; // c7t317i31
	assign leaf[442] = !f[677] && !f[595] && f[542] && f[241]; // c7t317i31
	assign leaf[443] = !f[677] && f[595] && !f[292] && !f[681]; // c7t317i31
	assign leaf[444] = !f[677] && f[595] && !f[292] && f[681]; // c7t317i31
	assign leaf[445] = !f[677] && f[595] && f[292]; // c7t317i31
	assign leaf[446] = f[677] && !f[682] && !f[516]; // c7t317i31
	assign leaf[447] = f[677] && !f[682] && f[516] && !f[234]; // c7t317i31
	assign leaf[448] = f[677] && !f[682] && f[516] && f[234]; // c7t317i31
	assign leaf[449] = f[677] && f[682]; // c7t317i31
	assign leaf[450] = !f[609] && !f[549] && !f[206] && !f[260]; // c7t327i32
	assign leaf[451] = !f[609] && !f[549] && !f[206] && f[260]; // c7t327i32
	assign leaf[452] = !f[609] && !f[549] && f[206] && !f[634]; // c7t327i32
	assign leaf[453] = !f[609] && !f[549] && f[206] && f[634]; // c7t327i32
	assign leaf[454] = !f[609] && f[549] && !f[434] && !f[626]; // c7t327i32
	assign leaf[455] = !f[609] && f[549] && !f[434] && f[626]; // c7t327i32
	assign leaf[456] = !f[609] && f[549] && f[434] && !f[202]; // c7t327i32
	assign leaf[457] = !f[609] && f[549] && f[434] && f[202]; // c7t327i32
	assign leaf[458] = f[609] && !f[319] && !f[720]; // c7t327i32
	assign leaf[459] = f[609] && !f[319] && f[720] && !f[294]; // c7t327i32
	assign leaf[460] = f[609] && !f[319] && f[720] && f[294]; // c7t327i32
	assign leaf[461] = f[609] && f[319] && !f[262]; // c7t327i32
	assign leaf[462] = f[609] && f[319] && f[262] && !f[397]; // c7t327i32
	assign leaf[463] = f[609] && f[319] && f[262] && f[397]; // c7t327i32
	assign leaf[464] = !f[242] && !f[411] && !f[177] && !f[231]; // c7t337i33
	assign leaf[465] = !f[242] && !f[411] && !f[177] && f[231]; // c7t337i33
	assign leaf[466] = !f[242] && !f[411] && f[177] && !f[492]; // c7t337i33
	assign leaf[467] = !f[242] && !f[411] && f[177] && f[492]; // c7t337i33
	assign leaf[468] = !f[242] && f[411] && !f[323] && !f[463]; // c7t337i33
	assign leaf[469] = !f[242] && f[411] && !f[323] && f[463]; // c7t337i33
	assign leaf[470] = !f[242] && f[411] && f[323] && !f[550]; // c7t337i33
	assign leaf[471] = !f[242] && f[411] && f[323] && f[550]; // c7t337i33
	assign leaf[472] = f[242] && !f[240] && !f[236] && !f[156]; // c7t337i33
	assign leaf[473] = f[242] && !f[240] && !f[236] && f[156]; // c7t337i33
	assign leaf[474] = f[242] && !f[240] && f[236] && !f[322]; // c7t337i33
	assign leaf[475] = f[242] && !f[240] && f[236] && f[322]; // c7t337i33
	assign leaf[476] = f[242] && f[240] && !f[349] && !f[325]; // c7t337i33
	assign leaf[477] = f[242] && f[240] && !f[349] && f[325]; // c7t337i33
	assign leaf[478] = f[242] && f[240] && f[349] && !f[267]; // c7t337i33
	assign leaf[479] = f[242] && f[240] && f[349] && f[267]; // c7t337i33
	assign leaf[480] = !f[460] && !f[515] && !f[379] && !f[569]; // c7t347i34
	assign leaf[481] = !f[460] && !f[515] && !f[379] && f[569]; // c7t347i34
	assign leaf[482] = !f[460] && !f[515] && f[379] && !f[349]; // c7t347i34
	assign leaf[483] = !f[460] && !f[515] && f[379] && f[349]; // c7t347i34
	assign leaf[484] = !f[460] && f[515] && !f[678] && !f[234]; // c7t347i34
	assign leaf[485] = !f[460] && f[515] && !f[678] && f[234]; // c7t347i34
	assign leaf[486] = !f[460] && f[515] && f[678] && !f[262]; // c7t347i34
	assign leaf[487] = !f[460] && f[515] && f[678] && f[262]; // c7t347i34
	assign leaf[488] = f[460] && !f[372] && !f[374] && !f[342]; // c7t347i34
	assign leaf[489] = f[460] && !f[372] && !f[374] && f[342]; // c7t347i34
	assign leaf[490] = f[460] && !f[372] && f[374] && !f[497]; // c7t347i34
	assign leaf[491] = f[460] && !f[372] && f[374] && f[497]; // c7t347i34
	assign leaf[492] = f[460] && f[372] && !f[471] && !f[568]; // c7t347i34
	assign leaf[493] = f[460] && f[372] && !f[471] && f[568]; // c7t347i34
	assign leaf[494] = f[460] && f[372] && f[471] && !f[549]; // c7t347i34
	assign leaf[495] = f[460] && f[372] && f[471] && f[549]; // c7t347i34
	assign leaf[496] = !f[555] && !f[129] && !f[635] && !f[437]; // c7t357i35
	assign leaf[497] = !f[555] && !f[129] && !f[635] && f[437]; // c7t357i35
	assign leaf[498] = !f[555] && !f[129] && f[635] && !f[319]; // c7t357i35
	assign leaf[499] = !f[555] && !f[129] && f[635] && f[319]; // c7t357i35
	assign leaf[500] = !f[555] && f[129]; // c7t357i35
	assign leaf[501] = f[555] && !f[540]; // c7t357i35
	assign leaf[502] = f[555] && f[540]; // c7t357i35
	assign leaf[503] = !f[127] && !f[677] && !f[595] && !f[515]; // c7t367i36
	assign leaf[504] = !f[127] && !f[677] && !f[595] && f[515]; // c7t367i36
	assign leaf[505] = !f[127] && !f[677] && f[595] && !f[406]; // c7t367i36
	assign leaf[506] = !f[127] && !f[677] && f[595] && f[406]; // c7t367i36
	assign leaf[507] = !f[127] && f[677] && !f[576] && !f[541]; // c7t367i36
	assign leaf[508] = !f[127] && f[677] && !f[576] && f[541]; // c7t367i36
	assign leaf[509] = !f[127] && f[677] && f[576]; // c7t367i36
	assign leaf[510] = f[127] && !f[539]; // c7t367i36
	assign leaf[511] = f[127] && f[539]; // c7t367i36
	assign leaf[512] = !f[256] && !f[663] && !f[349] && !f[433]; // c7t377i37
	assign leaf[513] = !f[256] && !f[663] && !f[349] && f[433]; // c7t377i37
	assign leaf[514] = !f[256] && !f[663] && f[349] && !f[384]; // c7t377i37
	assign leaf[515] = !f[256] && !f[663] && f[349] && f[384]; // c7t377i37
	assign leaf[516] = !f[256] && f[663] && !f[263] && !f[178]; // c7t377i37
	assign leaf[517] = !f[256] && f[663] && !f[263] && f[178]; // c7t377i37
	assign leaf[518] = !f[256] && f[663] && f[263] && !f[489]; // c7t377i37
	assign leaf[519] = !f[256] && f[663] && f[263] && f[489]; // c7t377i37
	assign leaf[520] = f[256] && !f[287] && !f[659] && !f[494]; // c7t377i37
	assign leaf[521] = f[256] && !f[287] && !f[659] && f[494]; // c7t377i37
	assign leaf[522] = f[256] && !f[287] && f[659]; // c7t377i37
	assign leaf[523] = f[256] && f[287] && !f[554] && !f[294]; // c7t377i37
	assign leaf[524] = f[256] && f[287] && !f[554] && f[294]; // c7t377i37
	assign leaf[525] = f[256] && f[287] && f[554]; // c7t377i37
	assign leaf[526] = !f[122] && !f[160] && !f[129] && !f[325]; // c7t387i38
	assign leaf[527] = !f[122] && !f[160] && !f[129] && f[325]; // c7t387i38
	assign leaf[528] = !f[122] && !f[160] && f[129]; // c7t387i38
	assign leaf[529] = !f[122] && f[160] && !f[684]; // c7t387i38
	assign leaf[530] = !f[122] && f[160] && f[684]; // c7t387i38
	assign leaf[531] = f[122]; // c7t387i38
	assign leaf[532] = !f[124] && !f[459] && !f[183] && !f[151]; // c7t397i39
	assign leaf[533] = !f[124] && !f[459] && !f[183] && f[151]; // c7t397i39
	assign leaf[534] = !f[124] && !f[459] && f[183] && !f[321]; // c7t397i39
	assign leaf[535] = !f[124] && !f[459] && f[183] && f[321]; // c7t397i39
	assign leaf[536] = !f[124] && f[459] && !f[400] && !f[324]; // c7t397i39
	assign leaf[537] = !f[124] && f[459] && !f[400] && f[324]; // c7t397i39
	assign leaf[538] = !f[124] && f[459] && f[400] && !f[469]; // c7t397i39
	assign leaf[539] = !f[124] && f[459] && f[400] && f[469]; // c7t397i39
	assign leaf[540] = f[124]; // c7t397i39
	assign leaf[541] = !f[510] && !f[411] && !f[242] && !f[467]; // c7t407i40
	assign leaf[542] = !f[510] && !f[411] && !f[242] && f[467]; // c7t407i40
	assign leaf[543] = !f[510] && !f[411] && f[242] && !f[578]; // c7t407i40
	assign leaf[544] = !f[510] && !f[411] && f[242] && f[578]; // c7t407i40
	assign leaf[545] = !f[510] && f[411] && !f[383] && !f[551]; // c7t407i40
	assign leaf[546] = !f[510] && f[411] && !f[383] && f[551]; // c7t407i40
	assign leaf[547] = !f[510] && f[411] && f[383] && !f[460]; // c7t407i40
	assign leaf[548] = !f[510] && f[411] && f[383] && f[460]; // c7t407i40
	assign leaf[549] = f[510] && !f[257] && !f[541] && !f[519]; // c7t407i40
	assign leaf[550] = f[510] && !f[257] && !f[541] && f[519]; // c7t407i40
	assign leaf[551] = f[510] && !f[257] && f[541] && !f[219]; // c7t407i40
	assign leaf[552] = f[510] && !f[257] && f[541] && f[219]; // c7t407i40
	assign leaf[553] = f[510] && f[257]; // c7t407i40
	assign leaf[554] = !f[158] && !f[637] && !f[202] && !f[549]; // c7t417i41
	assign leaf[555] = !f[158] && !f[637] && !f[202] && f[549]; // c7t417i41
	assign leaf[556] = !f[158] && !f[637] && f[202] && !f[493]; // c7t417i41
	assign leaf[557] = !f[158] && !f[637] && f[202] && f[493]; // c7t417i41
	assign leaf[558] = !f[158] && f[637] && !f[318]; // c7t417i41
	assign leaf[559] = !f[158] && f[637] && f[318] && !f[179]; // c7t417i41
	assign leaf[560] = !f[158] && f[637] && f[318] && f[179]; // c7t417i41
	assign leaf[561] = f[158] && !f[154] && !f[232] && !f[377]; // c7t417i41
	assign leaf[562] = f[158] && !f[154] && !f[232] && f[377]; // c7t417i41
	assign leaf[563] = f[158] && !f[154] && f[232]; // c7t417i41
	assign leaf[564] = f[158] && f[154] && !f[235]; // c7t417i41
	assign leaf[565] = f[158] && f[154] && f[235] && !f[263]; // c7t417i41
	assign leaf[566] = f[158] && f[154] && f[235] && f[263]; // c7t417i41
	assign leaf[567] = !f[677] && !f[595] && !f[434] && !f[378]; // c7t427i42
	assign leaf[568] = !f[677] && !f[595] && !f[434] && f[378]; // c7t427i42
	assign leaf[569] = !f[677] && !f[595] && f[434] && !f[351]; // c7t427i42
	assign leaf[570] = !f[677] && !f[595] && f[434] && f[351]; // c7t427i42
	assign leaf[571] = !f[677] && f[595] && !f[573] && !f[656]; // c7t427i42
	assign leaf[572] = !f[677] && f[595] && !f[573] && f[656]; // c7t427i42
	assign leaf[573] = !f[677] && f[595] && f[573]; // c7t427i42
	assign leaf[574] = f[677] && !f[404] && !f[681] && !f[234]; // c7t427i42
	assign leaf[575] = f[677] && !f[404] && !f[681] && f[234]; // c7t427i42
	assign leaf[576] = f[677] && !f[404] && f[681]; // c7t427i42
	assign leaf[577] = f[677] && f[404]; // c7t427i42
	assign leaf[578] = !f[438] && !f[214] && !f[301] && !f[349]; // c7t437i43
	assign leaf[579] = !f[438] && !f[214] && !f[301] && f[349]; // c7t437i43
	assign leaf[580] = !f[438] && !f[214] && f[301] && !f[541]; // c7t437i43
	assign leaf[581] = !f[438] && !f[214] && f[301] && f[541]; // c7t437i43
	assign leaf[582] = !f[438] && f[214] && !f[544] && !f[681]; // c7t437i43
	assign leaf[583] = !f[438] && f[214] && !f[544] && f[681]; // c7t437i43
	assign leaf[584] = !f[438] && f[214] && f[544] && !f[152]; // c7t437i43
	assign leaf[585] = !f[438] && f[214] && f[544] && f[152]; // c7t437i43
	assign leaf[586] = f[438] && !f[202] && !f[515] && !f[596]; // c7t437i43
	assign leaf[587] = f[438] && !f[202] && !f[515] && f[596]; // c7t437i43
	assign leaf[588] = f[438] && !f[202] && f[515] && !f[318]; // c7t437i43
	assign leaf[589] = f[438] && !f[202] && f[515] && f[318]; // c7t437i43
	assign leaf[590] = f[438] && f[202] && !f[257] && !f[598]; // c7t437i43
	assign leaf[591] = f[438] && f[202] && !f[257] && f[598]; // c7t437i43
	assign leaf[592] = f[438] && f[202] && f[257] && !f[260]; // c7t437i43
	assign leaf[593] = f[438] && f[202] && f[257] && f[260]; // c7t437i43
	assign leaf[594] = !f[715] && !f[576] && !f[632] && !f[179]; // c7t447i44
	assign leaf[595] = !f[715] && !f[576] && !f[632] && f[179]; // c7t447i44
	assign leaf[596] = !f[715] && !f[576] && f[632] && !f[716]; // c7t447i44
	assign leaf[597] = !f[715] && !f[576] && f[632] && f[716]; // c7t447i44
	assign leaf[598] = !f[715] && f[576] && !f[230] && !f[406]; // c7t447i44
	assign leaf[599] = !f[715] && f[576] && !f[230] && f[406]; // c7t447i44
	assign leaf[600] = !f[715] && f[576] && f[230] && !f[492]; // c7t447i44
	assign leaf[601] = !f[715] && f[576] && f[230] && f[492]; // c7t447i44
	assign leaf[602] = f[715] && !f[631] && !f[181] && !f[518]; // c7t447i44
	assign leaf[603] = f[715] && !f[631] && !f[181] && f[518]; // c7t447i44
	assign leaf[604] = f[715] && !f[631] && f[181] && !f[322]; // c7t447i44
	assign leaf[605] = f[715] && !f[631] && f[181] && f[322]; // c7t447i44
	assign leaf[606] = f[715] && f[631] && !f[518] && !f[436]; // c7t447i44
	assign leaf[607] = f[715] && f[631] && !f[518] && f[436]; // c7t447i44
	assign leaf[608] = f[715] && f[631] && f[518] && !f[302]; // c7t447i44
	assign leaf[609] = f[715] && f[631] && f[518] && f[302]; // c7t447i44
	assign leaf[610] = !f[128] && !f[241] && !f[322] && !f[434]; // c7t457i45
	assign leaf[611] = !f[128] && !f[241] && !f[322] && f[434]; // c7t457i45
	assign leaf[612] = !f[128] && !f[241] && f[322] && !f[412]; // c7t457i45
	assign leaf[613] = !f[128] && !f[241] && f[322] && f[412]; // c7t457i45
	assign leaf[614] = !f[128] && f[241] && !f[239] && !f[154]; // c7t457i45
	assign leaf[615] = !f[128] && f[241] && !f[239] && f[154]; // c7t457i45
	assign leaf[616] = !f[128] && f[241] && f[239] && !f[207]; // c7t457i45
	assign leaf[617] = !f[128] && f[241] && f[239] && f[207]; // c7t457i45
	assign leaf[618] = f[128]; // c7t457i45
	assign leaf[619] = !f[256] && !f[663] && !f[177] && !f[232]; // c7t467i46
	assign leaf[620] = !f[256] && !f[663] && !f[177] && f[232]; // c7t467i46
	assign leaf[621] = !f[256] && !f[663] && f[177] && !f[183]; // c7t467i46
	assign leaf[622] = !f[256] && !f[663] && f[177] && f[183]; // c7t467i46
	assign leaf[623] = !f[256] && f[663] && !f[263] && !f[550]; // c7t467i46
	assign leaf[624] = !f[256] && f[663] && !f[263] && f[550]; // c7t467i46
	assign leaf[625] = !f[256] && f[663] && f[263] && !f[459]; // c7t467i46
	assign leaf[626] = !f[256] && f[663] && f[263] && f[459]; // c7t467i46
	assign leaf[627] = f[256] && !f[493] && !f[436]; // c7t467i46
	assign leaf[628] = f[256] && !f[493] && f[436] && !f[239]; // c7t467i46
	assign leaf[629] = f[256] && !f[493] && f[436] && f[239]; // c7t467i46
	assign leaf[630] = f[256] && f[493] && !f[581] && !f[552]; // c7t467i46
	assign leaf[631] = f[256] && f[493] && !f[581] && f[552]; // c7t467i46
	assign leaf[632] = f[256] && f[493] && f[581]; // c7t467i46
	assign leaf[633] = !f[295] && !f[350] && !f[213] && !f[435]; // c7t477i47
	assign leaf[634] = !f[295] && !f[350] && !f[213] && f[435]; // c7t477i47
	assign leaf[635] = !f[295] && !f[350] && f[213] && !f[461]; // c7t477i47
	assign leaf[636] = !f[295] && !f[350] && f[213] && f[461]; // c7t477i47
	assign leaf[637] = !f[295] && f[350] && !f[210] && !f[266]; // c7t477i47
	assign leaf[638] = !f[295] && f[350] && !f[210] && f[266]; // c7t477i47
	assign leaf[639] = !f[295] && f[350] && f[210] && !f[460]; // c7t477i47
	assign leaf[640] = !f[295] && f[350] && f[210] && f[460]; // c7t477i47
	assign leaf[641] = f[295] && !f[404] && !f[491] && !f[212]; // c7t477i47
	assign leaf[642] = f[295] && !f[404] && !f[491] && f[212]; // c7t477i47
	assign leaf[643] = f[295] && !f[404] && f[491] && !f[658]; // c7t477i47
	assign leaf[644] = f[295] && !f[404] && f[491] && f[658]; // c7t477i47
	assign leaf[645] = f[295] && f[404] && !f[345] && !f[569]; // c7t477i47
	assign leaf[646] = f[295] && f[404] && !f[345] && f[569]; // c7t477i47
	assign leaf[647] = f[295] && f[404] && f[345] && !f[406]; // c7t477i47
	assign leaf[648] = f[295] && f[404] && f[345] && f[406]; // c7t477i47
	assign leaf[649] = !f[128] && !f[296] && !f[431] && !f[485]; // c7t487i48
	assign leaf[650] = !f[128] && !f[296] && !f[431] && f[485]; // c7t487i48
	assign leaf[651] = !f[128] && !f[296] && f[431] && !f[457]; // c7t487i48
	assign leaf[652] = !f[128] && !f[296] && f[431] && f[457]; // c7t487i48
	assign leaf[653] = !f[128] && f[296] && !f[404] && !f[492]; // c7t487i48
	assign leaf[654] = !f[128] && f[296] && !f[404] && f[492]; // c7t487i48
	assign leaf[655] = !f[128] && f[296] && f[404] && !f[318]; // c7t487i48
	assign leaf[656] = !f[128] && f[296] && f[404] && f[318]; // c7t487i48
	assign leaf[657] = f[128]; // c7t487i48
	assign leaf[658] = !f[125] && !f[244] && !f[527] && !f[324]; // c7t497i49
	assign leaf[659] = !f[125] && !f[244] && !f[527] && f[324]; // c7t497i49
	assign leaf[660] = !f[125] && !f[244] && f[527] && !f[404]; // c7t497i49
	assign leaf[661] = !f[125] && !f[244] && f[527] && f[404]; // c7t497i49
	assign leaf[662] = !f[125] && f[244] && !f[604] && !f[207]; // c7t497i49
	assign leaf[663] = !f[125] && f[244] && !f[604] && f[207]; // c7t497i49
	assign leaf[664] = !f[125] && f[244] && f[604] && !f[494]; // c7t497i49
	assign leaf[665] = !f[125] && f[244] && f[604] && f[494]; // c7t497i49
	assign leaf[666] = f[125] && !f[486]; // c7t497i49
	assign leaf[667] = f[125] && f[486]; // c7t497i49
	assign leaf[668] = !f[743] && !f[354] && !f[239] && !f[358]; // c7t507i50
	assign leaf[669] = !f[743] && !f[354] && !f[239] && f[358]; // c7t507i50
	assign leaf[670] = !f[743] && !f[354] && f[239] && !f[549]; // c7t507i50
	assign leaf[671] = !f[743] && !f[354] && f[239] && f[549]; // c7t507i50
	assign leaf[672] = !f[743] && f[354] && !f[459] && !f[401]; // c7t507i50
	assign leaf[673] = !f[743] && f[354] && !f[459] && f[401]; // c7t507i50
	assign leaf[674] = !f[743] && f[354] && f[459] && !f[401]; // c7t507i50
	assign leaf[675] = !f[743] && f[354] && f[459] && f[401]; // c7t507i50
	assign leaf[676] = f[743] && !f[264] && !f[231] && !f[716]; // c7t507i50
	assign leaf[677] = f[743] && !f[264] && !f[231] && f[716]; // c7t507i50
	assign leaf[678] = f[743] && !f[264] && f[231]; // c7t507i50
	assign leaf[679] = f[743] && f[264] && !f[343] && !f[235]; // c7t507i50
	assign leaf[680] = f[743] && f[264] && !f[343] && f[235]; // c7t507i50
	assign leaf[681] = f[743] && f[264] && f[343] && !f[260]; // c7t507i50
	assign leaf[682] = f[743] && f[264] && f[343] && f[260]; // c7t507i50
	assign leaf[683] = !f[690] && !f[634] && !f[177] && !f[232]; // c7t517i51
	assign leaf[684] = !f[690] && !f[634] && !f[177] && f[232]; // c7t517i51
	assign leaf[685] = !f[690] && !f[634] && f[177] && !f[523]; // c7t517i51
	assign leaf[686] = !f[690] && !f[634] && f[177] && f[523]; // c7t517i51
	assign leaf[687] = !f[690] && f[634] && !f[434] && !f[342]; // c7t517i51
	assign leaf[688] = !f[690] && f[634] && !f[434] && f[342]; // c7t517i51
	assign leaf[689] = !f[690] && f[634] && f[434] && !f[468]; // c7t517i51
	assign leaf[690] = !f[690] && f[634] && f[434] && f[468]; // c7t517i51
	assign leaf[691] = f[690] && !f[291] && !f[522] && !f[633]; // c7t517i51
	assign leaf[692] = f[690] && !f[291] && !f[522] && f[633]; // c7t517i51
	assign leaf[693] = f[690] && !f[291] && f[522] && !f[496]; // c7t517i51
	assign leaf[694] = f[690] && !f[291] && f[522] && f[496]; // c7t517i51
	assign leaf[695] = f[690] && f[291] && !f[489] && !f[686]; // c7t517i51
	assign leaf[696] = f[690] && f[291] && !f[489] && f[686]; // c7t517i51
	assign leaf[697] = f[690] && f[291] && f[489] && !f[286]; // c7t517i51
	assign leaf[698] = f[690] && f[291] && f[489] && f[286]; // c7t517i51
	assign leaf[699] = !f[242] && !f[457] && !f[397] && !f[347]; // c7t527i52
	assign leaf[700] = !f[242] && !f[457] && !f[397] && f[347]; // c7t527i52
	assign leaf[701] = !f[242] && !f[457] && f[397] && !f[513]; // c7t527i52
	assign leaf[702] = !f[242] && !f[457] && f[397] && f[513]; // c7t527i52
	assign leaf[703] = !f[242] && f[457] && !f[399] && !f[322]; // c7t527i52
	assign leaf[704] = !f[242] && f[457] && !f[399] && f[322]; // c7t527i52
	assign leaf[705] = !f[242] && f[457] && f[399] && !f[347]; // c7t527i52
	assign leaf[706] = !f[242] && f[457] && f[399] && f[347]; // c7t527i52
	assign leaf[707] = f[242] && !f[604] && !f[320] && !f[317]; // c7t527i52
	assign leaf[708] = f[242] && !f[604] && !f[320] && f[317]; // c7t527i52
	assign leaf[709] = f[242] && !f[604] && f[320] && !f[373]; // c7t527i52
	assign leaf[710] = f[242] && !f[604] && f[320] && f[373]; // c7t527i52
	assign leaf[711] = f[242] && f[604] && !f[716] && !f[655]; // c7t527i52
	assign leaf[712] = f[242] && f[604] && !f[716] && f[655]; // c7t527i52
	assign leaf[713] = f[242] && f[604] && f[716] && !f[515]; // c7t527i52
	assign leaf[714] = f[242] && f[604] && f[716] && f[515]; // c7t527i52
	assign leaf[715] = !f[160] && !f[639] && !f[528] && !f[434]; // c7t537i53
	assign leaf[716] = !f[160] && !f[639] && !f[528] && f[434]; // c7t537i53
	assign leaf[717] = !f[160] && !f[639] && f[528] && !f[381]; // c7t537i53
	assign leaf[718] = !f[160] && !f[639] && f[528] && f[381]; // c7t537i53
	assign leaf[719] = !f[160] && f[639]; // c7t537i53
	assign leaf[720] = f[160] && !f[182]; // c7t537i53
	assign leaf[721] = f[160] && f[182]; // c7t537i53
	assign leaf[722] = !f[678] && !f[596] && !f[434] && !f[488]; // c7t547i54
	assign leaf[723] = !f[678] && !f[596] && !f[434] && f[488]; // c7t547i54
	assign leaf[724] = !f[678] && !f[596] && f[434] && !f[490]; // c7t547i54
	assign leaf[725] = !f[678] && !f[596] && f[434] && f[490]; // c7t547i54
	assign leaf[726] = !f[678] && f[596] && !f[542] && !f[399]; // c7t547i54
	assign leaf[727] = !f[678] && f[596] && !f[542] && f[399]; // c7t547i54
	assign leaf[728] = !f[678] && f[596] && f[542] && !f[546]; // c7t547i54
	assign leaf[729] = !f[678] && f[596] && f[542] && f[546]; // c7t547i54
	assign leaf[730] = f[678] && !f[597] && !f[325]; // c7t547i54
	assign leaf[731] = f[678] && !f[597] && f[325]; // c7t547i54
	assign leaf[732] = f[678] && f[597] && !f[521] && !f[404]; // c7t547i54
	assign leaf[733] = f[678] && f[597] && !f[521] && f[404]; // c7t547i54
	assign leaf[734] = f[678] && f[597] && f[521]; // c7t547i54
	assign leaf[735] = !f[122] && !f[148] && !f[160] && !f[600]; // c7t557i55
	assign leaf[736] = !f[122] && !f[148] && !f[160] && f[600]; // c7t557i55
	assign leaf[737] = !f[122] && !f[148] && f[160] && !f[651]; // c7t557i55
	assign leaf[738] = !f[122] && !f[148] && f[160] && f[651]; // c7t557i55
	assign leaf[739] = !f[122] && f[148] && !f[153] && !f[173]; // c7t557i55
	assign leaf[740] = !f[122] && f[148] && !f[153] && f[173]; // c7t557i55
	assign leaf[741] = !f[122] && f[148] && f[153] && !f[548]; // c7t557i55
	assign leaf[742] = !f[122] && f[148] && f[153] && f[548]; // c7t557i55
	assign leaf[743] = f[122]; // c7t557i55
	assign leaf[744] = !f[583] && !f[122] && !f[183] && !f[488]; // c7t567i56
	assign leaf[745] = !f[583] && !f[122] && !f[183] && f[488]; // c7t567i56
	assign leaf[746] = !f[583] && !f[122] && f[183] && !f[320]; // c7t567i56
	assign leaf[747] = !f[583] && !f[122] && f[183] && f[320]; // c7t567i56
	assign leaf[748] = !f[583] && f[122]; // c7t567i56
	assign leaf[749] = f[583]; // c7t567i56
	assign leaf[750] = !f[359] && !f[202] && !f[548] && !f[603]; // c7t577i57
	assign leaf[751] = !f[359] && !f[202] && !f[548] && f[603]; // c7t577i57
	assign leaf[752] = !f[359] && !f[202] && f[548] && !f[433]; // c7t577i57
	assign leaf[753] = !f[359] && !f[202] && f[548] && f[433]; // c7t577i57
	assign leaf[754] = !f[359] && f[202] && !f[492] && !f[205]; // c7t577i57
	assign leaf[755] = !f[359] && f[202] && !f[492] && f[205]; // c7t577i57
	assign leaf[756] = !f[359] && f[202] && f[492] && !f[540]; // c7t577i57
	assign leaf[757] = !f[359] && f[202] && f[492] && f[540]; // c7t577i57
	assign leaf[758] = f[359] && !f[240] && !f[542] && !f[319]; // c7t577i57
	assign leaf[759] = f[359] && !f[240] && !f[542] && f[319]; // c7t577i57
	assign leaf[760] = f[359] && !f[240] && f[542]; // c7t577i57
	assign leaf[761] = f[359] && f[240] && !f[466] && !f[545]; // c7t577i57
	assign leaf[762] = f[359] && f[240] && !f[466] && f[545]; // c7t577i57
	assign leaf[763] = f[359] && f[240] && f[466] && !f[710]; // c7t577i57
	assign leaf[764] = f[359] && f[240] && f[466] && f[710]; // c7t577i57
	assign leaf[765] = !f[191] && !f[126] && !f[608] && !f[295]; // c7t587i58
	assign leaf[766] = !f[191] && !f[126] && !f[608] && f[295]; // c7t587i58
	assign leaf[767] = !f[191] && !f[126] && f[608] && !f[270]; // c7t587i58
	assign leaf[768] = !f[191] && !f[126] && f[608] && f[270]; // c7t587i58
	assign leaf[769] = !f[191] && f[126] && !f[629]; // c7t587i58
	assign leaf[770] = !f[191] && f[126] && f[629]; // c7t587i58
	assign leaf[771] = f[191] && !f[679]; // c7t587i58
	assign leaf[772] = f[191] && f[679]; // c7t587i58
	assign leaf[773] = !f[129] && !f[122] && !f[432] && !f[377]; // c7t597i59
	assign leaf[774] = !f[129] && !f[122] && !f[432] && f[377]; // c7t597i59
	assign leaf[775] = !f[129] && !f[122] && f[432] && !f[345]; // c7t597i59
	assign leaf[776] = !f[129] && !f[122] && f[432] && f[345]; // c7t597i59
	assign leaf[777] = !f[129] && f[122]; // c7t597i59
	assign leaf[778] = f[129]; // c7t597i59
	assign leaf[779] = !f[239] && !f[236] && !f[327] && !f[156]; // c7t607i60
	assign leaf[780] = !f[239] && !f[236] && !f[327] && f[156]; // c7t607i60
	assign leaf[781] = !f[239] && !f[236] && f[327] && !f[206]; // c7t607i60
	assign leaf[782] = !f[239] && !f[236] && f[327] && f[206]; // c7t607i60
	assign leaf[783] = !f[239] && f[236] && !f[247] && !f[685]; // c7t607i60
	assign leaf[784] = !f[239] && f[236] && !f[247] && f[685]; // c7t607i60
	assign leaf[785] = !f[239] && f[236] && f[247]; // c7t607i60
	assign leaf[786] = f[239] && !f[371] && !f[369] && !f[457]; // c7t607i60
	assign leaf[787] = f[239] && !f[371] && !f[369] && f[457]; // c7t607i60
	assign leaf[788] = f[239] && !f[371] && f[369] && !f[489]; // c7t607i60
	assign leaf[789] = f[239] && !f[371] && f[369] && f[489]; // c7t607i60
	assign leaf[790] = f[239] && f[371] && !f[460] && !f[293]; // c7t607i60
	assign leaf[791] = f[239] && f[371] && !f[460] && f[293]; // c7t607i60
	assign leaf[792] = f[239] && f[371] && f[460] && !f[428]; // c7t607i60
	assign leaf[793] = f[239] && f[371] && f[460] && f[428]; // c7t607i60
	assign leaf[794] = !f[582] && !f[161] && !f[272] && !f[355]; // c7t617i61
	assign leaf[795] = !f[582] && !f[161] && !f[272] && f[355]; // c7t617i61
	assign leaf[796] = !f[582] && !f[161] && f[272] && !f[406]; // c7t617i61
	assign leaf[797] = !f[582] && !f[161] && f[272] && f[406]; // c7t617i61
	assign leaf[798] = !f[582] && f[161]; // c7t617i61
	assign leaf[799] = f[582] && !f[350] && !f[212]; // c7t617i61
	assign leaf[800] = f[582] && !f[350] && f[212]; // c7t617i61
	assign leaf[801] = f[582] && f[350]; // c7t617i61
	assign leaf[802] = !f[638] && !f[348] && !f[374] && !f[185]; // c7t627i62
	assign leaf[803] = !f[638] && !f[348] && !f[374] && f[185]; // c7t627i62
	assign leaf[804] = !f[638] && !f[348] && f[374] && !f[460]; // c7t627i62
	assign leaf[805] = !f[638] && !f[348] && f[374] && f[460]; // c7t627i62
	assign leaf[806] = !f[638] && f[348] && !f[401] && !f[210]; // c7t627i62
	assign leaf[807] = !f[638] && f[348] && !f[401] && f[210]; // c7t627i62
	assign leaf[808] = !f[638] && f[348] && f[401] && !f[460]; // c7t627i62
	assign leaf[809] = !f[638] && f[348] && f[401] && f[460]; // c7t627i62
	assign leaf[810] = f[638]; // c7t627i62
	assign leaf[811] = !f[372] && !f[405] && !f[492] && !f[205]; // c7t637i63
	assign leaf[812] = !f[372] && !f[405] && !f[492] && f[205]; // c7t637i63
	assign leaf[813] = !f[372] && !f[405] && f[492] && !f[398]; // c7t637i63
	assign leaf[814] = !f[372] && !f[405] && f[492] && f[398]; // c7t637i63
	assign leaf[815] = !f[372] && f[405] && !f[346] && !f[435]; // c7t637i63
	assign leaf[816] = !f[372] && f[405] && !f[346] && f[435]; // c7t637i63
	assign leaf[817] = !f[372] && f[405] && f[346] && !f[316]; // c7t637i63
	assign leaf[818] = !f[372] && f[405] && f[346] && f[316]; // c7t637i63
	assign leaf[819] = f[372] && !f[460] && !f[318] && !f[349]; // c7t637i63
	assign leaf[820] = f[372] && !f[460] && !f[318] && f[349]; // c7t637i63
	assign leaf[821] = f[372] && !f[460] && f[318] && !f[516]; // c7t637i63
	assign leaf[822] = f[372] && !f[460] && f[318] && f[516]; // c7t637i63
	assign leaf[823] = f[372] && f[460] && !f[470] && !f[458]; // c7t637i63
	assign leaf[824] = f[372] && f[460] && !f[470] && f[458]; // c7t637i63
	assign leaf[825] = f[372] && f[460] && f[470] && !f[577]; // c7t637i63
	assign leaf[826] = f[372] && f[460] && f[470] && f[577]; // c7t637i63
	assign leaf[827] = !f[325] && !f[205] && !f[542] && !f[314]; // c7t647i64
	assign leaf[828] = !f[325] && !f[205] && !f[542] && f[314]; // c7t647i64
	assign leaf[829] = !f[325] && !f[205] && f[542] && !f[677]; // c7t647i64
	assign leaf[830] = !f[325] && !f[205] && f[542] && f[677]; // c7t647i64
	assign leaf[831] = !f[325] && f[205] && !f[605] && !f[575]; // c7t647i64
	assign leaf[832] = !f[325] && f[205] && !f[605] && f[575]; // c7t647i64
	assign leaf[833] = !f[325] && f[205] && f[605] && !f[263]; // c7t647i64
	assign leaf[834] = !f[325] && f[205] && f[605] && f[263]; // c7t647i64
	assign leaf[835] = f[325] && !f[150] && !f[437] && !f[548]; // c7t647i64
	assign leaf[836] = f[325] && !f[150] && !f[437] && f[548]; // c7t647i64
	assign leaf[837] = f[325] && !f[150] && f[437] && !f[176]; // c7t647i64
	assign leaf[838] = f[325] && !f[150] && f[437] && f[176]; // c7t647i64
	assign leaf[839] = f[325] && f[150] && !f[233] && !f[463]; // c7t647i64
	assign leaf[840] = f[325] && f[150] && !f[233] && f[463]; // c7t647i64
	assign leaf[841] = f[325] && f[150] && f[233] && !f[430]; // c7t647i64
	assign leaf[842] = f[325] && f[150] && f[233] && f[430]; // c7t647i64
	assign leaf[843] = !f[269] && !f[601] && !f[684] && !f[545]; // c7t657i65
	assign leaf[844] = !f[269] && !f[601] && !f[684] && f[545]; // c7t657i65
	assign leaf[845] = !f[269] && !f[601] && f[684] && !f[660]; // c7t657i65
	assign leaf[846] = !f[269] && !f[601] && f[684] && f[660]; // c7t657i65
	assign leaf[847] = !f[269] && f[601] && !f[177] && !f[453]; // c7t657i65
	assign leaf[848] = !f[269] && f[601] && !f[177] && f[453]; // c7t657i65
	assign leaf[849] = !f[269] && f[601] && f[177] && !f[550]; // c7t657i65
	assign leaf[850] = !f[269] && f[601] && f[177] && f[550]; // c7t657i65
	assign leaf[851] = f[269] && !f[577] && !f[663] && !f[482]; // c7t657i65
	assign leaf[852] = f[269] && !f[577] && !f[663] && f[482]; // c7t657i65
	assign leaf[853] = f[269] && !f[577] && f[663] && !f[291]; // c7t657i65
	assign leaf[854] = f[269] && !f[577] && f[663] && f[291]; // c7t657i65
	assign leaf[855] = f[269] && f[577] && !f[522] && !f[465]; // c7t657i65
	assign leaf[856] = f[269] && f[577] && !f[522] && f[465]; // c7t657i65
	assign leaf[857] = f[269] && f[577] && f[522] && !f[660]; // c7t657i65
	assign leaf[858] = f[269] && f[577] && f[522] && f[660]; // c7t657i65
	assign leaf[859] = !f[129] && !f[148] && !f[160] && !f[150]; // c7t667i66
	assign leaf[860] = !f[129] && !f[148] && !f[160] && f[150]; // c7t667i66
	assign leaf[861] = !f[129] && !f[148] && f[160]; // c7t667i66
	assign leaf[862] = !f[129] && f[148] && !f[153] && !f[146]; // c7t667i66
	assign leaf[863] = !f[129] && f[148] && !f[153] && f[146]; // c7t667i66
	assign leaf[864] = !f[129] && f[148] && f[153] && !f[520]; // c7t667i66
	assign leaf[865] = !f[129] && f[148] && f[153] && f[520]; // c7t667i66
	assign leaf[866] = f[129]; // c7t667i66
	assign leaf[867] = !f[473] && !f[441] && !f[206] && !f[432]; // c7t677i67
	assign leaf[868] = !f[473] && !f[441] && !f[206] && f[432]; // c7t677i67
	assign leaf[869] = !f[473] && !f[441] && f[206] && !f[260]; // c7t677i67
	assign leaf[870] = !f[473] && !f[441] && f[206] && f[260]; // c7t677i67
	assign leaf[871] = !f[473] && f[441] && !f[542] && !f[241]; // c7t677i67
	assign leaf[872] = !f[473] && f[441] && !f[542] && f[241]; // c7t677i67
	assign leaf[873] = !f[473] && f[441] && f[542] && !f[651]; // c7t677i67
	assign leaf[874] = !f[473] && f[441] && f[542] && f[651]; // c7t677i67
	assign leaf[875] = f[473]; // c7t677i67
	assign leaf[876] = !f[528] && !f[510] && !f[527] && !f[274]; // c7t687i68
	assign leaf[877] = !f[528] && !f[510] && !f[527] && f[274]; // c7t687i68
	assign leaf[878] = !f[528] && !f[510] && f[527] && !f[242]; // c7t687i68
	assign leaf[879] = !f[528] && !f[510] && f[527] && f[242]; // c7t687i68
	assign leaf[880] = !f[528] && f[510] && !f[660] && !f[656]; // c7t687i68
	assign leaf[881] = !f[528] && f[510] && !f[660] && f[656]; // c7t687i68
	assign leaf[882] = !f[528] && f[510] && f[660] && !f[457]; // c7t687i68
	assign leaf[883] = !f[528] && f[510] && f[660] && f[457]; // c7t687i68
	assign leaf[884] = f[528] && !f[353]; // c7t687i68
	assign leaf[885] = f[528] && f[353]; // c7t687i68
	assign leaf[886] = !f[269] && !f[519] && !f[210] && !f[318]; // c7t697i69
	assign leaf[887] = !f[269] && !f[519] && !f[210] && f[318]; // c7t697i69
	assign leaf[888] = !f[269] && !f[519] && f[210] && !f[373]; // c7t697i69
	assign leaf[889] = !f[269] && !f[519] && f[210] && f[373]; // c7t697i69
	assign leaf[890] = !f[269] && f[519] && !f[205] && !f[324]; // c7t697i69
	assign leaf[891] = !f[269] && f[519] && !f[205] && f[324]; // c7t697i69
	assign leaf[892] = !f[269] && f[519] && f[205] && !f[211]; // c7t697i69
	assign leaf[893] = !f[269] && f[519] && f[205] && f[211]; // c7t697i69
	assign leaf[894] = f[269] && !f[173] && !f[349] && !f[370]; // c7t697i69
	assign leaf[895] = f[269] && !f[173] && !f[349] && f[370]; // c7t697i69
	assign leaf[896] = f[269] && !f[173] && f[349] && !f[266]; // c7t697i69
	assign leaf[897] = f[269] && !f[173] && f[349] && f[266]; // c7t697i69
	assign leaf[898] = f[269] && f[173] && !f[550]; // c7t697i69
	assign leaf[899] = f[269] && f[173] && f[550]; // c7t697i69
	assign leaf[900] = !f[214] && !f[543] && !f[457] && !f[370]; // c7t707i70
	assign leaf[901] = !f[214] && !f[543] && !f[457] && f[370]; // c7t707i70
	assign leaf[902] = !f[214] && !f[543] && f[457] && !f[488]; // c7t707i70
	assign leaf[903] = !f[214] && !f[543] && f[457] && f[488]; // c7t707i70
	assign leaf[904] = !f[214] && f[543] && !f[679] && !f[528]; // c7t707i70
	assign leaf[905] = !f[214] && f[543] && !f[679] && f[528]; // c7t707i70
	assign leaf[906] = !f[214] && f[543] && f[679]; // c7t707i70
	assign leaf[907] = f[214] && !f[577] && !f[269] && !f[323]; // c7t707i70
	assign leaf[908] = f[214] && !f[577] && !f[269] && f[323]; // c7t707i70
	assign leaf[909] = f[214] && !f[577] && f[269] && !f[236]; // c7t707i70
	assign leaf[910] = f[214] && !f[577] && f[269] && f[236]; // c7t707i70
	assign leaf[911] = f[214] && f[577] && !f[716] && !f[715]; // c7t707i70
	assign leaf[912] = f[214] && f[577] && !f[716] && f[715]; // c7t707i70
	assign leaf[913] = f[214] && f[577] && f[716] && !f[261]; // c7t707i70
	assign leaf[914] = f[214] && f[577] && f[716] && f[261]; // c7t707i70
	assign leaf[915] = !f[494] && !f[605] && !f[690] && !f[575]; // c7t717i71
	assign leaf[916] = !f[494] && !f[605] && !f[690] && f[575]; // c7t717i71
	assign leaf[917] = !f[494] && !f[605] && f[690] && !f[440]; // c7t717i71
	assign leaf[918] = !f[494] && !f[605] && f[690] && f[440]; // c7t717i71
	assign leaf[919] = !f[494] && f[605] && !f[285] && !f[455]; // c7t717i71
	assign leaf[920] = !f[494] && f[605] && !f[285] && f[455]; // c7t717i71
	assign leaf[921] = !f[494] && f[605] && f[285] && !f[579]; // c7t717i71
	assign leaf[922] = !f[494] && f[605] && f[285] && f[579]; // c7t717i71
	assign leaf[923] = f[494] && !f[571] && !f[655] && !f[576]; // c7t717i71
	assign leaf[924] = f[494] && !f[571] && !f[655] && f[576]; // c7t717i71
	assign leaf[925] = f[494] && !f[571] && f[655] && !f[518]; // c7t717i71
	assign leaf[926] = f[494] && !f[571] && f[655] && f[518]; // c7t717i71
	assign leaf[927] = f[494] && f[571] && !f[654] && !f[173]; // c7t717i71
	assign leaf[928] = f[494] && f[571] && !f[654] && f[173]; // c7t717i71
	assign leaf[929] = f[494] && f[571] && f[654] && !f[516]; // c7t717i71
	assign leaf[930] = f[494] && f[571] && f[654] && f[516]; // c7t717i71
	assign leaf[931] = !f[359] && !f[663] && !f[320] && !f[317]; // c7t727i72
	assign leaf[932] = !f[359] && !f[663] && !f[320] && f[317]; // c7t727i72
	assign leaf[933] = !f[359] && !f[663] && f[320] && !f[318]; // c7t727i72
	assign leaf[934] = !f[359] && !f[663] && f[320] && f[318]; // c7t727i72
	assign leaf[935] = !f[359] && f[663] && !f[577] && !f[178]; // c7t727i72
	assign leaf[936] = !f[359] && f[663] && !f[577] && f[178]; // c7t727i72
	assign leaf[937] = !f[359] && f[663] && f[577] && !f[516]; // c7t727i72
	assign leaf[938] = !f[359] && f[663] && f[577] && f[516]; // c7t727i72
	assign leaf[939] = f[359] && !f[456] && !f[369]; // c7t727i72
	assign leaf[940] = f[359] && !f[456] && f[369]; // c7t727i72
	assign leaf[941] = f[359] && f[456] && !f[485]; // c7t727i72
	assign leaf[942] = f[359] && f[456] && f[485]; // c7t727i72
	assign leaf[943] = !f[154] && !f[159] && !f[461] && !f[378]; // c7t737i73
	assign leaf[944] = !f[154] && !f[159] && !f[461] && f[378]; // c7t737i73
	assign leaf[945] = !f[154] && !f[159] && f[461] && !f[378]; // c7t737i73
	assign leaf[946] = !f[154] && !f[159] && f[461] && f[378]; // c7t737i73
	assign leaf[947] = !f[154] && f[159] && !f[263]; // c7t737i73
	assign leaf[948] = !f[154] && f[159] && f[263]; // c7t737i73
	assign leaf[949] = f[154] && !f[236] && !f[262] && !f[260]; // c7t737i73
	assign leaf[950] = f[154] && !f[236] && !f[262] && f[260]; // c7t737i73
	assign leaf[951] = f[154] && !f[236] && f[262]; // c7t737i73
	assign leaf[952] = f[154] && f[236] && !f[684] && !f[232]; // c7t737i73
	assign leaf[953] = f[154] && f[236] && !f[684] && f[232]; // c7t737i73
	assign leaf[954] = f[154] && f[236] && f[684] && !f[234]; // c7t737i73
	assign leaf[955] = f[154] && f[236] && f[684] && f[234]; // c7t737i73
	assign leaf[956] = !f[709] && !f[129] && !f[214] && !f[323]; // c7t747i74
	assign leaf[957] = !f[709] && !f[129] && !f[214] && f[323]; // c7t747i74
	assign leaf[958] = !f[709] && !f[129] && f[214] && !f[320]; // c7t747i74
	assign leaf[959] = !f[709] && !f[129] && f[214] && f[320]; // c7t747i74
	assign leaf[960] = !f[709] && f[129]; // c7t747i74
	assign leaf[961] = f[709] && !f[654] && !f[271]; // c7t747i74
	assign leaf[962] = f[709] && !f[654] && f[271]; // c7t747i74
	assign leaf[963] = f[709] && f[654] && !f[322] && !f[303]; // c7t747i74
	assign leaf[964] = f[709] && f[654] && !f[322] && f[303]; // c7t747i74
	assign leaf[965] = f[709] && f[654] && f[322] && !f[329]; // c7t747i74
	assign leaf[966] = f[709] && f[654] && f[322] && f[329]; // c7t747i74
	assign leaf[967] = !f[515] && !f[457] && !f[426] && !f[265]; // c7t757i75
	assign leaf[968] = !f[515] && !f[457] && !f[426] && f[265]; // c7t757i75
	assign leaf[969] = !f[515] && !f[457] && f[426] && !f[430]; // c7t757i75
	assign leaf[970] = !f[515] && !f[457] && f[426] && f[430]; // c7t757i75
	assign leaf[971] = !f[515] && f[457] && !f[460] && !f[569]; // c7t757i75
	assign leaf[972] = !f[515] && f[457] && !f[460] && f[569]; // c7t757i75
	assign leaf[973] = !f[515] && f[457] && f[460] && !f[372]; // c7t757i75
	assign leaf[974] = !f[515] && f[457] && f[460] && f[372]; // c7t757i75
	assign leaf[975] = f[515] && !f[428] && !f[426] && !f[291]; // c7t757i75
	assign leaf[976] = f[515] && !f[428] && !f[426] && f[291]; // c7t757i75
	assign leaf[977] = f[515] && !f[428] && f[426]; // c7t757i75
	assign leaf[978] = f[515] && f[428] && !f[485] && !f[601]; // c7t757i75
	assign leaf[979] = f[515] && f[428] && !f[485] && f[601]; // c7t757i75
	assign leaf[980] = f[515] && f[428] && f[485] && !f[405]; // c7t757i75
	assign leaf[981] = f[515] && f[428] && f[485] && f[405]; // c7t757i75
	assign leaf[982] = !f[510] && !f[464] && !f[547] && !f[176]; // c7t767i76
	assign leaf[983] = !f[510] && !f[464] && !f[547] && f[176]; // c7t767i76
	assign leaf[984] = !f[510] && !f[464] && f[547] && !f[377]; // c7t767i76
	assign leaf[985] = !f[510] && !f[464] && f[547] && f[377]; // c7t767i76
	assign leaf[986] = !f[510] && f[464] && !f[383] && !f[518]; // c7t767i76
	assign leaf[987] = !f[510] && f[464] && !f[383] && f[518]; // c7t767i76
	assign leaf[988] = !f[510] && f[464] && f[383] && !f[326]; // c7t767i76
	assign leaf[989] = !f[510] && f[464] && f[383] && f[326]; // c7t767i76
	assign leaf[990] = f[510] && !f[685] && !f[661] && !f[314]; // c7t767i76
	assign leaf[991] = f[510] && !f[685] && !f[661] && f[314]; // c7t767i76
	assign leaf[992] = f[510] && !f[685] && f[661]; // c7t767i76
	assign leaf[993] = f[510] && f[685] && !f[296]; // c7t767i76
	assign leaf[994] = f[510] && f[685] && f[296]; // c7t767i76
	assign leaf[995] = !f[528] && !f[527] && !f[709] && !f[708]; // c7t777i77
	assign leaf[996] = !f[528] && !f[527] && !f[709] && f[708]; // c7t777i77
	assign leaf[997] = !f[528] && !f[527] && f[709] && !f[630]; // c7t777i77
	assign leaf[998] = !f[528] && !f[527] && f[709] && f[630]; // c7t777i77
	assign leaf[999] = !f[528] && f[527] && !f[242]; // c7t777i77
	assign leaf[1000] = !f[528] && f[527] && f[242]; // c7t777i77
	assign leaf[1001] = f[528] && !f[600]; // c7t777i77
	assign leaf[1002] = f[528] && f[600]; // c7t777i77
	assign leaf[1003] = !f[452] && !f[577] && !f[689] && !f[180]; // c7t787i78
	assign leaf[1004] = !f[452] && !f[577] && !f[689] && f[180]; // c7t787i78
	assign leaf[1005] = !f[452] && !f[577] && f[689] && !f[686]; // c7t787i78
	assign leaf[1006] = !f[452] && !f[577] && f[689] && f[686]; // c7t787i78
	assign leaf[1007] = !f[452] && f[577] && !f[626] && !f[202]; // c7t787i78
	assign leaf[1008] = !f[452] && f[577] && !f[626] && f[202]; // c7t787i78
	assign leaf[1009] = !f[452] && f[577] && f[626] && !f[157]; // c7t787i78
	assign leaf[1010] = !f[452] && f[577] && f[626] && f[157]; // c7t787i78
	assign leaf[1011] = f[452] && !f[427]; // c7t787i78
	assign leaf[1012] = f[452] && f[427]; // c7t787i78
	assign leaf[1013] = !f[437] && !f[273] && !f[176] && !f[517]; // c7t797i79
	assign leaf[1014] = !f[437] && !f[273] && !f[176] && f[517]; // c7t797i79
	assign leaf[1015] = !f[437] && !f[273] && f[176] && !f[494]; // c7t797i79
	assign leaf[1016] = !f[437] && !f[273] && f[176] && f[494]; // c7t797i79
	assign leaf[1017] = !f[437] && f[273] && !f[485] && !f[183]; // c7t797i79
	assign leaf[1018] = !f[437] && f[273] && !f[485] && f[183]; // c7t797i79
	assign leaf[1019] = !f[437] && f[273] && f[485]; // c7t797i79
	assign leaf[1020] = f[437] && !f[581] && !f[359] && !f[184]; // c7t797i79
	assign leaf[1021] = f[437] && !f[581] && !f[359] && f[184]; // c7t797i79
	assign leaf[1022] = f[437] && !f[581] && f[359] && !f[325]; // c7t797i79
	assign leaf[1023] = f[437] && !f[581] && f[359] && f[325]; // c7t797i79
	assign leaf[1024] = f[437] && f[581] && !f[204]; // c7t797i79
	assign leaf[1025] = f[437] && f[581] && f[204]; // c7t797i79
	assign leaf[1026] = !f[148] && !f[569] && !f[554] && !f[434]; // c7t807i80
	assign leaf[1027] = !f[148] && !f[569] && !f[554] && f[434]; // c7t807i80
	assign leaf[1028] = !f[148] && !f[569] && f[554] && !f[212]; // c7t807i80
	assign leaf[1029] = !f[148] && !f[569] && f[554] && f[212]; // c7t807i80
	assign leaf[1030] = !f[148] && f[569] && !f[651] && !f[260]; // c7t807i80
	assign leaf[1031] = !f[148] && f[569] && !f[651] && f[260]; // c7t807i80
	assign leaf[1032] = !f[148] && f[569] && f[651] && !f[547]; // c7t807i80
	assign leaf[1033] = !f[148] && f[569] && f[651] && f[547]; // c7t807i80
	assign leaf[1034] = f[148] && !f[324]; // c7t807i80
	assign leaf[1035] = f[148] && f[324] && !f[292] && !f[522]; // c7t807i80
	assign leaf[1036] = f[148] && f[324] && !f[292] && f[522]; // c7t807i80
	assign leaf[1037] = f[148] && f[324] && f[292]; // c7t807i80
	assign leaf[1038] = !f[154] && !f[266] && !f[575] && !f[269]; // c7t817i81
	assign leaf[1039] = !f[154] && !f[266] && !f[575] && f[269]; // c7t817i81
	assign leaf[1040] = !f[154] && !f[266] && f[575] && !f[205]; // c7t817i81
	assign leaf[1041] = !f[154] && !f[266] && f[575] && f[205]; // c7t817i81
	assign leaf[1042] = !f[154] && f[266] && !f[263] && !f[294]; // c7t817i81
	assign leaf[1043] = !f[154] && f[266] && !f[263] && f[294]; // c7t817i81
	assign leaf[1044] = !f[154] && f[266] && f[263] && !f[368]; // c7t817i81
	assign leaf[1045] = !f[154] && f[266] && f[263] && f[368]; // c7t817i81
	assign leaf[1046] = f[154] && !f[463] && !f[571]; // c7t817i81
	assign leaf[1047] = f[154] && !f[463] && f[571]; // c7t817i81
	assign leaf[1048] = f[154] && f[463] && !f[403] && !f[236]; // c7t817i81
	assign leaf[1049] = f[154] && f[463] && !f[403] && f[236]; // c7t817i81
	assign leaf[1050] = f[154] && f[463] && f[403] && !f[152]; // c7t817i81
	assign leaf[1051] = f[154] && f[463] && f[403] && f[152]; // c7t817i81
	assign leaf[1052] = !f[686] && !f[575] && !f[683] && !f[518]; // c7t827i82
	assign leaf[1053] = !f[686] && !f[575] && !f[683] && f[518]; // c7t827i82
	assign leaf[1054] = !f[686] && !f[575] && f[683] && !f[624]; // c7t827i82
	assign leaf[1055] = !f[686] && !f[575] && f[683] && f[624]; // c7t827i82
	assign leaf[1056] = !f[686] && f[575] && !f[492] && !f[203]; // c7t827i82
	assign leaf[1057] = !f[686] && f[575] && !f[492] && f[203]; // c7t827i82
	assign leaf[1058] = !f[686] && f[575] && f[492] && !f[259]; // c7t827i82
	assign leaf[1059] = !f[686] && f[575] && f[492] && f[259]; // c7t827i82
	assign leaf[1060] = f[686] && !f[682] && !f[661] && !f[323]; // c7t827i82
	assign leaf[1061] = f[686] && !f[682] && !f[661] && f[323]; // c7t827i82
	assign leaf[1062] = f[686] && !f[682] && f[661] && !f[716]; // c7t827i82
	assign leaf[1063] = f[686] && !f[682] && f[661] && f[716]; // c7t827i82
	assign leaf[1064] = f[686] && f[682] && !f[301] && !f[573]; // c7t827i82
	assign leaf[1065] = f[686] && f[682] && !f[301] && f[573]; // c7t827i82
	assign leaf[1066] = f[686] && f[682] && f[301]; // c7t827i82
	assign leaf[1067] = !f[238] && !f[235] && !f[322] && !f[208]; // c7t837i83
	assign leaf[1068] = !f[238] && !f[235] && !f[322] && f[208]; // c7t837i83
	assign leaf[1069] = !f[238] && !f[235] && f[322] && !f[318]; // c7t837i83
	assign leaf[1070] = !f[238] && !f[235] && f[322] && f[318]; // c7t837i83
	assign leaf[1071] = !f[238] && f[235] && !f[208] && !f[436]; // c7t837i83
	assign leaf[1072] = !f[238] && f[235] && !f[208] && f[436]; // c7t837i83
	assign leaf[1073] = !f[238] && f[235] && f[208] && !f[546]; // c7t837i83
	assign leaf[1074] = !f[238] && f[235] && f[208] && f[546]; // c7t837i83
	assign leaf[1075] = f[238] && !f[236] && !f[718] && !f[401]; // c7t837i83
	assign leaf[1076] = f[238] && !f[236] && !f[718] && f[401]; // c7t837i83
	assign leaf[1077] = f[238] && !f[236] && f[718]; // c7t837i83
	assign leaf[1078] = f[238] && f[236] && !f[329] && !f[214]; // c7t837i83
	assign leaf[1079] = f[238] && f[236] && !f[329] && f[214]; // c7t837i83
	assign leaf[1080] = f[238] && f[236] && f[329] && !f[274]; // c7t837i83
	assign leaf[1081] = f[238] && f[236] && f[329] && f[274]; // c7t837i83
	assign leaf[1082] = !f[464] && !f[574] && !f[300] && !f[236]; // c7t847i84
	assign leaf[1083] = !f[464] && !f[574] && !f[300] && f[236]; // c7t847i84
	assign leaf[1084] = !f[464] && !f[574] && f[300] && !f[683]; // c7t847i84
	assign leaf[1085] = !f[464] && !f[574] && f[300] && f[683]; // c7t847i84
	assign leaf[1086] = !f[464] && f[574] && !f[377] && !f[492]; // c7t847i84
	assign leaf[1087] = !f[464] && f[574] && !f[377] && f[492]; // c7t847i84
	assign leaf[1088] = !f[464] && f[574] && f[377] && !f[659]; // c7t847i84
	assign leaf[1089] = !f[464] && f[574] && f[377] && f[659]; // c7t847i84
	assign leaf[1090] = f[464] && !f[595] && !f[518] && !f[682]; // c7t847i84
	assign leaf[1091] = f[464] && !f[595] && !f[518] && f[682]; // c7t847i84
	assign leaf[1092] = f[464] && !f[595] && f[518] && !f[269]; // c7t847i84
	assign leaf[1093] = f[464] && !f[595] && f[518] && f[269]; // c7t847i84
	assign leaf[1094] = f[464] && f[595] && !f[677] && !f[440]; // c7t847i84
	assign leaf[1095] = f[464] && f[595] && !f[677] && f[440]; // c7t847i84
	assign leaf[1096] = f[464] && f[595] && f[677]; // c7t847i84
	assign leaf[1097] = !f[510] && !f[609] && !f[291] && !f[288]; // c7t857i85
	assign leaf[1098] = !f[510] && !f[609] && !f[291] && f[288]; // c7t857i85
	assign leaf[1099] = !f[510] && !f[609] && f[291] && !f[287]; // c7t857i85
	assign leaf[1100] = !f[510] && !f[609] && f[291] && f[287]; // c7t857i85
	assign leaf[1101] = !f[510] && f[609] && !f[349]; // c7t857i85
	assign leaf[1102] = !f[510] && f[609] && f[349]; // c7t857i85
	assign leaf[1103] = f[510] && !f[685] && !f[342] && !f[267]; // c7t857i85
	assign leaf[1104] = f[510] && !f[685] && !f[342] && f[267]; // c7t857i85
	assign leaf[1105] = f[510] && !f[685] && f[342]; // c7t857i85
	assign leaf[1106] = f[510] && f[685]; // c7t857i85
	assign leaf[1107] = !f[707] && !f[625] && !f[600] && !f[682]; // c7t867i86
	assign leaf[1108] = !f[707] && !f[625] && !f[600] && f[682]; // c7t867i86
	assign leaf[1109] = !f[707] && !f[625] && f[600] && !f[318]; // c7t867i86
	assign leaf[1110] = !f[707] && !f[625] && f[600] && f[318]; // c7t867i86
	assign leaf[1111] = !f[707] && f[625] && !f[602] && !f[685]; // c7t867i86
	assign leaf[1112] = !f[707] && f[625] && !f[602] && f[685]; // c7t867i86
	assign leaf[1113] = !f[707] && f[625] && f[602] && !f[685]; // c7t867i86
	assign leaf[1114] = !f[707] && f[625] && f[602] && f[685]; // c7t867i86
	assign leaf[1115] = f[707] && !f[597] && !f[706] && !f[185]; // c7t867i86
	assign leaf[1116] = f[707] && !f[597] && !f[706] && f[185]; // c7t867i86
	assign leaf[1117] = f[707] && !f[597] && f[706]; // c7t867i86
	assign leaf[1118] = f[707] && f[597] && !f[348] && !f[318]; // c7t867i86
	assign leaf[1119] = f[707] && f[597] && !f[348] && f[318]; // c7t867i86
	assign leaf[1120] = f[707] && f[597] && f[348]; // c7t867i86
	assign leaf[1121] = !f[434] && !f[488] && !f[458] && !f[432]; // c7t877i87
	assign leaf[1122] = !f[434] && !f[488] && !f[458] && f[432]; // c7t877i87
	assign leaf[1123] = !f[434] && !f[488] && f[458] && !f[374]; // c7t877i87
	assign leaf[1124] = !f[434] && !f[488] && f[458] && f[374]; // c7t877i87
	assign leaf[1125] = !f[434] && f[488] && !f[430] && !f[412]; // c7t877i87
	assign leaf[1126] = !f[434] && f[488] && !f[430] && f[412]; // c7t877i87
	assign leaf[1127] = !f[434] && f[488] && f[430] && !f[494]; // c7t877i87
	assign leaf[1128] = !f[434] && f[488] && f[430] && f[494]; // c7t877i87
	assign leaf[1129] = f[434] && !f[606] && !f[320] && !f[346]; // c7t877i87
	assign leaf[1130] = f[434] && !f[606] && !f[320] && f[346]; // c7t877i87
	assign leaf[1131] = f[434] && !f[606] && f[320] && !f[210]; // c7t877i87
	assign leaf[1132] = f[434] && !f[606] && f[320] && f[210]; // c7t877i87
	assign leaf[1133] = f[434] && f[606] && !f[202]; // c7t877i87
	assign leaf[1134] = f[434] && f[606] && f[202] && !f[327]; // c7t877i87
	assign leaf[1135] = f[434] && f[606] && f[202] && f[327]; // c7t877i87
	assign leaf[1136] = !f[148] && !f[494] && !f[690] && !f[206]; // c7t887i88
	assign leaf[1137] = !f[148] && !f[494] && !f[690] && f[206]; // c7t887i88
	assign leaf[1138] = !f[148] && !f[494] && f[690] && !f[182]; // c7t887i88
	assign leaf[1139] = !f[148] && !f[494] && f[690] && f[182]; // c7t887i88
	assign leaf[1140] = !f[148] && f[494] && !f[346] && !f[185]; // c7t887i88
	assign leaf[1141] = !f[148] && f[494] && !f[346] && f[185]; // c7t887i88
	assign leaf[1142] = !f[148] && f[494] && f[346] && !f[407]; // c7t887i88
	assign leaf[1143] = !f[148] && f[494] && f[346] && f[407]; // c7t887i88
	assign leaf[1144] = f[148] && !f[356] && !f[211]; // c7t887i88
	assign leaf[1145] = f[148] && !f[356] && f[211] && !f[545]; // c7t887i88
	assign leaf[1146] = f[148] && !f[356] && f[211] && f[545]; // c7t887i88
	assign leaf[1147] = f[148] && f[356]; // c7t887i88
	assign leaf[1148] = !f[510] && !f[428] && !f[457] && !f[544]; // c7t897i89
	assign leaf[1149] = !f[510] && !f[428] && !f[457] && f[544]; // c7t897i89
	assign leaf[1150] = !f[510] && !f[428] && f[457] && !f[401]; // c7t897i89
	assign leaf[1151] = !f[510] && !f[428] && f[457] && f[401]; // c7t897i89
	assign leaf[1152] = !f[510] && f[428] && !f[515] && !f[460]; // c7t897i89
	assign leaf[1153] = !f[510] && f[428] && !f[515] && f[460]; // c7t897i89
	assign leaf[1154] = !f[510] && f[428] && f[515] && !f[468]; // c7t897i89
	assign leaf[1155] = !f[510] && f[428] && f[515] && f[468]; // c7t897i89
	assign leaf[1156] = f[510] && !f[685] && !f[342]; // c7t897i89
	assign leaf[1157] = f[510] && !f[685] && f[342]; // c7t897i89
	assign leaf[1158] = f[510] && f[685]; // c7t897i89
	assign leaf[1159] = !f[704] && !f[595] && !f[720] && !f[206]; // c7t907i90
	assign leaf[1160] = !f[704] && !f[595] && !f[720] && f[206]; // c7t907i90
	assign leaf[1161] = !f[704] && !f[595] && f[720] && !f[266]; // c7t907i90
	assign leaf[1162] = !f[704] && !f[595] && f[720] && f[266]; // c7t907i90
	assign leaf[1163] = !f[704] && f[595] && !f[573] && !f[434]; // c7t907i90
	assign leaf[1164] = !f[704] && f[595] && !f[573] && f[434]; // c7t907i90
	assign leaf[1165] = !f[704] && f[595] && f[573] && !f[294]; // c7t907i90
	assign leaf[1166] = !f[704] && f[595] && f[573] && f[294]; // c7t907i90
	assign leaf[1167] = f[704]; // c7t907i90
	assign leaf[1168] = !f[148] && !f[312] && !f[463] && !f[601]; // c7t917i91
	assign leaf[1169] = !f[148] && !f[312] && !f[463] && f[601]; // c7t917i91
	assign leaf[1170] = !f[148] && !f[312] && f[463] && !f[578]; // c7t917i91
	assign leaf[1171] = !f[148] && !f[312] && f[463] && f[578]; // c7t917i91
	assign leaf[1172] = !f[148] && f[312] && !f[553] && !f[398]; // c7t917i91
	assign leaf[1173] = !f[148] && f[312] && !f[553] && f[398]; // c7t917i91
	assign leaf[1174] = !f[148] && f[312] && f[553]; // c7t917i91
	assign leaf[1175] = f[148] && !f[630] && !f[184]; // c7t917i91
	assign leaf[1176] = f[148] && !f[630] && f[184]; // c7t917i91
	assign leaf[1177] = f[148] && f[630] && !f[655]; // c7t917i91
	assign leaf[1178] = f[148] && f[630] && f[655]; // c7t917i91
	assign leaf[1179] = !f[298] && !f[323] && !f[287] && !f[715]; // c7t927i92
	assign leaf[1180] = !f[298] && !f[323] && !f[287] && f[715]; // c7t927i92
	assign leaf[1181] = !f[298] && !f[323] && f[287] && !f[461]; // c7t927i92
	assign leaf[1182] = !f[298] && !f[323] && f[287] && f[461]; // c7t927i92
	assign leaf[1183] = !f[298] && f[323] && !f[687] && !f[431]; // c7t927i92
	assign leaf[1184] = !f[298] && f[323] && !f[687] && f[431]; // c7t927i92
	assign leaf[1185] = !f[298] && f[323] && f[687] && !f[347]; // c7t927i92
	assign leaf[1186] = !f[298] && f[323] && f[687] && f[347]; // c7t927i92
	assign leaf[1187] = f[298] && !f[406] && !f[158] && !f[351]; // c7t927i92
	assign leaf[1188] = f[298] && !f[406] && !f[158] && f[351]; // c7t927i92
	assign leaf[1189] = f[298] && !f[406] && f[158]; // c7t927i92
	assign leaf[1190] = f[298] && f[406] && !f[570] && !f[202]; // c7t927i92
	assign leaf[1191] = f[298] && f[406] && !f[570] && f[202]; // c7t927i92
	assign leaf[1192] = f[298] && f[406] && f[570] && !f[602]; // c7t927i92
	assign leaf[1193] = f[298] && f[406] && f[570] && f[602]; // c7t927i92
	assign leaf[1194] = !f[349] && !f[432] && !f[488] && !f[290]; // c7t937i93
	assign leaf[1195] = !f[349] && !f[432] && !f[488] && f[290]; // c7t937i93
	assign leaf[1196] = !f[349] && !f[432] && f[488] && !f[429]; // c7t937i93
	assign leaf[1197] = !f[349] && !f[432] && f[488] && f[429]; // c7t937i93
	assign leaf[1198] = !f[349] && f[432] && !f[319] && !f[463]; // c7t937i93
	assign leaf[1199] = !f[349] && f[432] && !f[319] && f[463]; // c7t937i93
	assign leaf[1200] = !f[349] && f[432] && f[319] && !f[286]; // c7t937i93
	assign leaf[1201] = !f[349] && f[432] && f[319] && f[286]; // c7t937i93
	assign leaf[1202] = f[349] && !f[234] && !f[264] && !f[570]; // c7t937i93
	assign leaf[1203] = f[349] && !f[234] && !f[264] && f[570]; // c7t937i93
	assign leaf[1204] = f[349] && !f[234] && f[264] && !f[430]; // c7t937i93
	assign leaf[1205] = f[349] && !f[234] && f[264] && f[430]; // c7t937i93
	assign leaf[1206] = f[349] && f[234] && !f[265] && !f[405]; // c7t937i93
	assign leaf[1207] = f[349] && f[234] && !f[265] && f[405]; // c7t937i93
	assign leaf[1208] = f[349] && f[234] && f[265] && !f[289]; // c7t937i93
	assign leaf[1209] = f[349] && f[234] && f[265] && f[289]; // c7t937i93
	assign leaf[1210] = !f[605] && !f[472] && !f[482] && !f[411]; // c7t947i94
	assign leaf[1211] = !f[605] && !f[472] && !f[482] && f[411]; // c7t947i94
	assign leaf[1212] = !f[605] && !f[472] && f[482] && !f[429]; // c7t947i94
	assign leaf[1213] = !f[605] && !f[472] && f[482] && f[429]; // c7t947i94
	assign leaf[1214] = !f[605] && f[472] && !f[431]; // c7t947i94
	assign leaf[1215] = !f[605] && f[472] && f[431]; // c7t947i94
	assign leaf[1216] = f[605] && !f[516] && !f[682] && !f[627]; // c7t947i94
	assign leaf[1217] = f[605] && !f[516] && !f[682] && f[627]; // c7t947i94
	assign leaf[1218] = f[605] && !f[516] && f[682]; // c7t947i94
	assign leaf[1219] = f[605] && f[516] && !f[524] && !f[216]; // c7t947i94
	assign leaf[1220] = f[605] && f[516] && !f[524] && f[216]; // c7t947i94
	assign leaf[1221] = f[605] && f[516] && f[524] && !f[688]; // c7t947i94
	assign leaf[1222] = f[605] && f[516] && f[524] && f[688]; // c7t947i94
	assign leaf[1223] = !f[241] && !f[350] && !f[434] && !f[349]; // c7t957i95
	assign leaf[1224] = !f[241] && !f[350] && !f[434] && f[349]; // c7t957i95
	assign leaf[1225] = !f[241] && !f[350] && f[434] && !f[653]; // c7t957i95
	assign leaf[1226] = !f[241] && !f[350] && f[434] && f[653]; // c7t957i95
	assign leaf[1227] = !f[241] && f[350] && !f[329] && !f[430]; // c7t957i95
	assign leaf[1228] = !f[241] && f[350] && !f[329] && f[430]; // c7t957i95
	assign leaf[1229] = !f[241] && f[350] && f[329] && !f[657]; // c7t957i95
	assign leaf[1230] = !f[241] && f[350] && f[329] && f[657]; // c7t957i95
	assign leaf[1231] = f[241] && !f[229] && !f[356] && !f[322]; // c7t957i95
	assign leaf[1232] = f[241] && !f[229] && !f[356] && f[322]; // c7t957i95
	assign leaf[1233] = f[241] && !f[229] && f[356] && !f[245]; // c7t957i95
	assign leaf[1234] = f[241] && !f[229] && f[356] && f[245]; // c7t957i95
	assign leaf[1235] = f[241] && f[229] && !f[541] && !f[627]; // c7t957i95
	assign leaf[1236] = f[241] && f[229] && !f[541] && f[627]; // c7t957i95
	assign leaf[1237] = f[241] && f[229] && f[541]; // c7t957i95
	assign leaf[1238] = !f[472] && !f[202] && !f[262] && !f[292]; // c7t967i96
	assign leaf[1239] = !f[472] && !f[202] && !f[262] && f[292]; // c7t967i96
	assign leaf[1240] = !f[472] && !f[202] && f[262] && !f[265]; // c7t967i96
	assign leaf[1241] = !f[472] && !f[202] && f[262] && f[265]; // c7t967i96
	assign leaf[1242] = !f[472] && f[202] && !f[568] && !f[598]; // c7t967i96
	assign leaf[1243] = !f[472] && f[202] && !f[568] && f[598]; // c7t967i96
	assign leaf[1244] = !f[472] && f[202] && f[568]; // c7t967i96
	assign leaf[1245] = f[472] && !f[457]; // c7t967i96
	assign leaf[1246] = f[472] && f[457]; // c7t967i96
	assign leaf[1247] = !f[359] && !f[206] && !f[260] && !f[154]; // c7t977i97
	assign leaf[1248] = !f[359] && !f[206] && !f[260] && f[154]; // c7t977i97
	assign leaf[1249] = !f[359] && !f[206] && f[260] && !f[291]; // c7t977i97
	assign leaf[1250] = !f[359] && !f[206] && f[260] && f[291]; // c7t977i97
	assign leaf[1251] = !f[359] && f[206] && !f[327] && !f[259]; // c7t977i97
	assign leaf[1252] = !f[359] && f[206] && !f[327] && f[259]; // c7t977i97
	assign leaf[1253] = !f[359] && f[206] && f[327] && !f[520]; // c7t977i97
	assign leaf[1254] = !f[359] && f[206] && f[327] && f[520]; // c7t977i97
	assign leaf[1255] = f[359] && !f[683] && !f[427]; // c7t977i97
	assign leaf[1256] = f[359] && !f[683] && f[427]; // c7t977i97
	assign leaf[1257] = f[359] && f[683]; // c7t977i97
	assign leaf[1258] = !f[154] && !f[159] && !f[182] && !f[542]; // c7t987i98
	assign leaf[1259] = !f[154] && !f[159] && !f[182] && f[542]; // c7t987i98
	assign leaf[1260] = !f[154] && !f[159] && f[182] && !f[290]; // c7t987i98
	assign leaf[1261] = !f[154] && !f[159] && f[182] && f[290]; // c7t987i98
	assign leaf[1262] = !f[154] && f[159]; // c7t987i98
	assign leaf[1263] = f[154] && !f[403] && !f[186] && !f[463]; // c7t987i98
	assign leaf[1264] = f[154] && !f[403] && !f[186] && f[463]; // c7t987i98
	assign leaf[1265] = f[154] && !f[403] && f[186] && !f[233]; // c7t987i98
	assign leaf[1266] = f[154] && !f[403] && f[186] && f[233]; // c7t987i98
	assign leaf[1267] = f[154] && f[403] && !f[684]; // c7t987i98
	assign leaf[1268] = f[154] && f[403] && f[684]; // c7t987i98
	assign leaf[1269] = !f[396] && !f[376] && !f[288] && !f[261]; // c7t997i99
	assign leaf[1270] = !f[396] && !f[376] && !f[288] && f[261]; // c7t997i99
	assign leaf[1271] = !f[396] && !f[376] && f[288] && !f[290]; // c7t997i99
	assign leaf[1272] = !f[396] && !f[376] && f[288] && f[290]; // c7t997i99
	assign leaf[1273] = !f[396] && f[376] && !f[289] && !f[402]; // c7t997i99
	assign leaf[1274] = !f[396] && f[376] && !f[289] && f[402]; // c7t997i99
	assign leaf[1275] = !f[396] && f[376] && f[289] && !f[293]; // c7t997i99
	assign leaf[1276] = !f[396] && f[376] && f[289] && f[293]; // c7t997i99
	assign leaf[1277] = f[396] && !f[346] && !f[491]; // c7t997i99
	assign leaf[1278] = f[396] && !f[346] && f[491]; // c7t997i99
	assign leaf[1279] = f[396] && f[346]; // c7t997i99
endmodule

module decision_tree_leaves_8(input logic [0:783] f, output logic [0:1497] leaf);
	assign leaf[0] = !f[487] && !f[488] && !f[486] && !f[489]; // c8t8i0
	assign leaf[1] = !f[487] && !f[488] && !f[486] && f[489]; // c8t8i0
	assign leaf[2] = !f[487] && !f[488] && f[486] && !f[377]; // c8t8i0
	assign leaf[3] = !f[487] && !f[488] && f[486] && f[377]; // c8t8i0
	assign leaf[4] = !f[487] && f[488] && !f[659] && !f[376]; // c8t8i0
	assign leaf[5] = !f[487] && f[488] && !f[659] && f[376]; // c8t8i0
	assign leaf[6] = !f[487] && f[488] && f[659] && !f[347]; // c8t8i0
	assign leaf[7] = !f[487] && f[488] && f[659] && f[347]; // c8t8i0
	assign leaf[8] = f[487] && !f[656] && !f[276] && !f[657]; // c8t8i0
	assign leaf[9] = f[487] && !f[656] && !f[276] && f[657]; // c8t8i0
	assign leaf[10] = f[487] && !f[656] && f[276] && !f[214]; // c8t8i0
	assign leaf[11] = f[487] && !f[656] && f[276] && f[214]; // c8t8i0
	assign leaf[12] = f[487] && f[656] && !f[405] && !f[457]; // c8t8i0
	assign leaf[13] = f[487] && f[656] && !f[405] && f[457]; // c8t8i0
	assign leaf[14] = f[487] && f[656] && f[405] && !f[514]; // c8t8i0
	assign leaf[15] = f[487] && f[656] && f[405] && f[514]; // c8t8i0
	assign leaf[16] = !f[376] && !f[349] && !f[403] && !f[276]; // c8t18i1
	assign leaf[17] = !f[376] && !f[349] && !f[403] && f[276]; // c8t18i1
	assign leaf[18] = !f[376] && !f[349] && f[403] && !f[515]; // c8t18i1
	assign leaf[19] = !f[376] && !f[349] && f[403] && f[515]; // c8t18i1
	assign leaf[20] = !f[376] && f[349] && !f[295] && !f[460]; // c8t18i1
	assign leaf[21] = !f[376] && f[349] && !f[295] && f[460]; // c8t18i1
	assign leaf[22] = !f[376] && f[349] && f[295] && !f[459]; // c8t18i1
	assign leaf[23] = !f[376] && f[349] && f[295] && f[459]; // c8t18i1
	assign leaf[24] = f[376] && !f[461] && !f[486] && !f[485]; // c8t18i1
	assign leaf[25] = f[376] && !f[461] && !f[486] && f[485]; // c8t18i1
	assign leaf[26] = f[376] && !f[461] && f[486] && !f[407]; // c8t18i1
	assign leaf[27] = f[376] && !f[461] && f[486] && f[407]; // c8t18i1
	assign leaf[28] = f[376] && f[461] && !f[657] && !f[623]; // c8t18i1
	assign leaf[29] = f[376] && f[461] && !f[657] && f[623]; // c8t18i1
	assign leaf[30] = f[376] && f[461] && f[657] && !f[515]; // c8t18i1
	assign leaf[31] = f[376] && f[461] && f[657] && f[515]; // c8t18i1
	assign leaf[32] = !f[657] && !f[275] && !f[376] && !f[629]; // c8t28i2
	assign leaf[33] = !f[657] && !f[275] && !f[376] && f[629]; // c8t28i2
	assign leaf[34] = !f[657] && !f[275] && f[376] && !f[662]; // c8t28i2
	assign leaf[35] = !f[657] && !f[275] && f[376] && f[662]; // c8t28i2
	assign leaf[36] = !f[657] && f[275] && !f[486] && !f[488]; // c8t28i2
	assign leaf[37] = !f[657] && f[275] && !f[486] && f[488]; // c8t28i2
	assign leaf[38] = !f[657] && f[275] && f[486] && !f[466]; // c8t28i2
	assign leaf[39] = !f[657] && f[275] && f[486] && f[466]; // c8t28i2
	assign leaf[40] = f[657] && !f[515] && !f[513] && !f[516]; // c8t28i2
	assign leaf[41] = f[657] && !f[515] && !f[513] && f[516]; // c8t28i2
	assign leaf[42] = f[657] && !f[515] && f[513] && !f[404]; // c8t28i2
	assign leaf[43] = f[657] && !f[515] && f[513] && f[404]; // c8t28i2
	assign leaf[44] = f[657] && f[515] && !f[433] && !f[378]; // c8t28i2
	assign leaf[45] = f[657] && f[515] && !f[433] && f[378]; // c8t28i2
	assign leaf[46] = f[657] && f[515] && f[433] && !f[573]; // c8t28i2
	assign leaf[47] = f[657] && f[515] && f[433] && f[573]; // c8t28i2
	assign leaf[48] = !f[405] && !f[432] && !f[378] && !f[460]; // c8t38i3
	assign leaf[49] = !f[405] && !f[432] && !f[378] && f[460]; // c8t38i3
	assign leaf[50] = !f[405] && !f[432] && f[378] && !f[488]; // c8t38i3
	assign leaf[51] = !f[405] && !f[432] && f[378] && f[488]; // c8t38i3
	assign leaf[52] = !f[405] && f[432] && !f[457] && !f[516]; // c8t38i3
	assign leaf[53] = !f[405] && f[432] && !f[457] && f[516]; // c8t38i3
	assign leaf[54] = !f[405] && f[432] && f[457] && !f[332]; // c8t38i3
	assign leaf[55] = !f[405] && f[432] && f[457] && f[332]; // c8t38i3
	assign leaf[56] = f[405] && !f[300] && !f[319] && !f[346]; // c8t38i3
	assign leaf[57] = f[405] && !f[300] && !f[319] && f[346]; // c8t38i3
	assign leaf[58] = f[405] && !f[300] && f[319] && !f[402]; // c8t38i3
	assign leaf[59] = f[405] && !f[300] && f[319] && f[402]; // c8t38i3
	assign leaf[60] = f[405] && f[300] && !f[438] && !f[183]; // c8t38i3
	assign leaf[61] = f[405] && f[300] && !f[438] && f[183]; // c8t38i3
	assign leaf[62] = f[405] && f[300] && f[438] && !f[660]; // c8t38i3
	assign leaf[63] = f[405] && f[300] && f[438] && f[660]; // c8t38i3
	assign leaf[64] = !f[433] && !f[431] && !f[434] && !f[429]; // c8t48i4
	assign leaf[65] = !f[433] && !f[431] && !f[434] && f[429]; // c8t48i4
	assign leaf[66] = !f[433] && !f[431] && f[434] && !f[377]; // c8t48i4
	assign leaf[67] = !f[433] && !f[431] && f[434] && f[377]; // c8t48i4
	assign leaf[68] = !f[433] && f[431] && !f[658] && !f[655]; // c8t48i4
	assign leaf[69] = !f[433] && f[431] && !f[658] && f[655]; // c8t48i4
	assign leaf[70] = !f[433] && f[431] && f[658] && !f[374]; // c8t48i4
	assign leaf[71] = !f[433] && f[431] && f[658] && f[374]; // c8t48i4
	assign leaf[72] = f[433] && !f[657] && !f[303] && !f[629]; // c8t48i4
	assign leaf[73] = f[433] && !f[657] && !f[303] && f[629]; // c8t48i4
	assign leaf[74] = f[433] && !f[657] && f[303] && !f[408]; // c8t48i4
	assign leaf[75] = f[433] && !f[657] && f[303] && f[408]; // c8t48i4
	assign leaf[76] = f[433] && f[657] && !f[515] && !f[512]; // c8t48i4
	assign leaf[77] = f[433] && f[657] && !f[515] && f[512]; // c8t48i4
	assign leaf[78] = f[433] && f[657] && f[515] && !f[290]; // c8t48i4
	assign leaf[79] = f[433] && f[657] && f[515] && f[290]; // c8t48i4
	assign leaf[80] = !f[433] && !f[431] && !f[378] && !f[405]; // c8t58i5
	assign leaf[81] = !f[433] && !f[431] && !f[378] && f[405]; // c8t58i5
	assign leaf[82] = !f[433] && !f[431] && f[378] && !f[489]; // c8t58i5
	assign leaf[83] = !f[433] && !f[431] && f[378] && f[489]; // c8t58i5
	assign leaf[84] = !f[433] && f[431] && !f[548] && !f[400]; // c8t58i5
	assign leaf[85] = !f[433] && f[431] && !f[548] && f[400]; // c8t58i5
	assign leaf[86] = !f[433] && f[431] && f[548] && !f[434]; // c8t58i5
	assign leaf[87] = !f[433] && f[431] && f[548] && f[434]; // c8t58i5
	assign leaf[88] = f[433] && !f[348] && !f[375] && !f[321]; // c8t58i5
	assign leaf[89] = f[433] && !f[348] && !f[375] && f[321]; // c8t58i5
	assign leaf[90] = f[433] && !f[348] && f[375] && !f[429]; // c8t58i5
	assign leaf[91] = f[433] && !f[348] && f[375] && f[429]; // c8t58i5
	assign leaf[92] = f[433] && f[348] && !f[402] && !f[294]; // c8t58i5
	assign leaf[93] = f[433] && f[348] && !f[402] && f[294]; // c8t58i5
	assign leaf[94] = f[433] && f[348] && f[402] && !f[289]; // c8t58i5
	assign leaf[95] = f[433] && f[348] && f[402] && f[289]; // c8t58i5
	assign leaf[96] = !f[406] && !f[404] && !f[430] && !f[350]; // c8t68i6
	assign leaf[97] = !f[406] && !f[404] && !f[430] && f[350]; // c8t68i6
	assign leaf[98] = !f[406] && !f[404] && f[430] && !f[493]; // c8t68i6
	assign leaf[99] = !f[406] && !f[404] && f[430] && f[493]; // c8t68i6
	assign leaf[100] = !f[406] && f[404] && !f[408] && !f[522]; // c8t68i6
	assign leaf[101] = !f[406] && f[404] && !f[408] && f[522]; // c8t68i6
	assign leaf[102] = !f[406] && f[404] && f[408] && !f[656]; // c8t68i6
	assign leaf[103] = !f[406] && f[404] && f[408] && f[656]; // c8t68i6
	assign leaf[104] = f[406] && !f[487] && !f[485] && !f[516]; // c8t68i6
	assign leaf[105] = f[406] && !f[487] && !f[485] && f[516]; // c8t68i6
	assign leaf[106] = f[406] && !f[487] && f[485] && !f[437]; // c8t68i6
	assign leaf[107] = f[406] && !f[487] && f[485] && f[437]; // c8t68i6
	assign leaf[108] = f[406] && f[487] && !f[428] && !f[348]; // c8t68i6
	assign leaf[109] = f[406] && f[487] && !f[428] && f[348]; // c8t68i6
	assign leaf[110] = f[406] && f[487] && f[428] && !f[625]; // c8t68i6
	assign leaf[111] = f[406] && f[487] && f[428] && f[625]; // c8t68i6
	assign leaf[112] = !f[658] && !f[652] && !f[686] && !f[303]; // c8t78i7
	assign leaf[113] = !f[658] && !f[652] && !f[686] && f[303]; // c8t78i7
	assign leaf[114] = !f[658] && !f[652] && f[686] && !f[571]; // c8t78i7
	assign leaf[115] = !f[658] && !f[652] && f[686] && f[571]; // c8t78i7
	assign leaf[116] = !f[658] && f[652] && !f[513] && !f[599]; // c8t78i7
	assign leaf[117] = !f[658] && f[652] && !f[513] && f[599]; // c8t78i7
	assign leaf[118] = !f[658] && f[652] && f[513] && !f[570]; // c8t78i7
	assign leaf[119] = !f[658] && f[652] && f[513] && f[570]; // c8t78i7
	assign leaf[120] = f[658] && !f[543] && !f[541] && !f[544]; // c8t78i7
	assign leaf[121] = f[658] && !f[543] && !f[541] && f[544]; // c8t78i7
	assign leaf[122] = f[658] && !f[543] && f[541] && !f[379]; // c8t78i7
	assign leaf[123] = f[658] && !f[543] && f[541] && f[379]; // c8t78i7
	assign leaf[124] = f[658] && f[543] && !f[484] && !f[601]; // c8t78i7
	assign leaf[125] = f[658] && f[543] && !f[484] && f[601]; // c8t78i7
	assign leaf[126] = f[658] && f[543] && f[484] && !f[303]; // c8t78i7
	assign leaf[127] = f[658] && f[543] && f[484] && f[303]; // c8t78i7
	assign leaf[128] = !f[439] && !f[267] && !f[349] && !f[375]; // c8t88i8
	assign leaf[129] = !f[439] && !f[267] && !f[349] && f[375]; // c8t88i8
	assign leaf[130] = !f[439] && !f[267] && f[349] && !f[406]; // c8t88i8
	assign leaf[131] = !f[439] && !f[267] && f[349] && f[406]; // c8t88i8
	assign leaf[132] = !f[439] && f[267] && !f[301] && !f[661]; // c8t88i8
	assign leaf[133] = !f[439] && f[267] && !f[301] && f[661]; // c8t88i8
	assign leaf[134] = !f[439] && f[267] && f[301] && !f[380]; // c8t88i8
	assign leaf[135] = !f[439] && f[267] && f[301] && f[380]; // c8t88i8
	assign leaf[136] = f[439] && !f[521] && !f[330] && !f[377]; // c8t88i8
	assign leaf[137] = f[439] && !f[521] && !f[330] && f[377]; // c8t88i8
	assign leaf[138] = f[439] && !f[521] && f[330] && !f[355]; // c8t88i8
	assign leaf[139] = f[439] && !f[521] && f[330] && f[355]; // c8t88i8
	assign leaf[140] = f[439] && f[521] && !f[304] && !f[154]; // c8t88i8
	assign leaf[141] = f[439] && f[521] && !f[304] && f[154]; // c8t88i8
	assign leaf[142] = f[439] && f[521] && f[304] && !f[468]; // c8t88i8
	assign leaf[143] = f[439] && f[521] && f[304] && f[468]; // c8t88i8
	assign leaf[144] = !f[658] && !f[624] && !f[686] && !f[630]; // c8t98i9
	assign leaf[145] = !f[658] && !f[624] && !f[686] && f[630]; // c8t98i9
	assign leaf[146] = !f[658] && !f[624] && f[686] && !f[516]; // c8t98i9
	assign leaf[147] = !f[658] && !f[624] && f[686] && f[516]; // c8t98i9
	assign leaf[148] = !f[658] && f[624] && !f[571] && !f[494]; // c8t98i9
	assign leaf[149] = !f[658] && f[624] && !f[571] && f[494]; // c8t98i9
	assign leaf[150] = !f[658] && f[624] && f[571] && !f[265]; // c8t98i9
	assign leaf[151] = !f[658] && f[624] && f[571] && f[265]; // c8t98i9
	assign leaf[152] = f[658] && !f[516] && !f[513] && !f[511]; // c8t98i9
	assign leaf[153] = f[658] && !f[516] && !f[513] && f[511]; // c8t98i9
	assign leaf[154] = f[658] && !f[516] && f[513] && !f[379]; // c8t98i9
	assign leaf[155] = f[658] && !f[516] && f[513] && f[379]; // c8t98i9
	assign leaf[156] = f[658] && f[516] && !f[602] && !f[514]; // c8t98i9
	assign leaf[157] = f[658] && f[516] && !f[602] && f[514]; // c8t98i9
	assign leaf[158] = f[658] && f[516] && f[602] && !f[317]; // c8t98i9
	assign leaf[159] = f[658] && f[516] && f[602] && f[317]; // c8t98i9
	assign leaf[160] = !f[439] && !f[302] && !f[183] && !f[154]; // c8t108i10
	assign leaf[161] = !f[439] && !f[302] && !f[183] && f[154]; // c8t108i10
	assign leaf[162] = !f[439] && !f[302] && f[183] && !f[299]; // c8t108i10
	assign leaf[163] = !f[439] && !f[302] && f[183] && f[299]; // c8t108i10
	assign leaf[164] = !f[439] && f[302] && !f[469] && !f[272]; // c8t108i10
	assign leaf[165] = !f[439] && f[302] && !f[469] && f[272]; // c8t108i10
	assign leaf[166] = !f[439] && f[302] && f[469] && !f[399]; // c8t108i10
	assign leaf[167] = !f[439] && f[302] && f[469] && f[399]; // c8t108i10
	assign leaf[168] = f[439] && !f[521] && !f[179] && !f[331]; // c8t108i10
	assign leaf[169] = f[439] && !f[521] && !f[179] && f[331]; // c8t108i10
	assign leaf[170] = f[439] && !f[521] && f[179] && !f[550]; // c8t108i10
	assign leaf[171] = f[439] && !f[521] && f[179] && f[550]; // c8t108i10
	assign leaf[172] = f[439] && f[521] && !f[304] && !f[378]; // c8t108i10
	assign leaf[173] = f[439] && f[521] && !f[304] && f[378]; // c8t108i10
	assign leaf[174] = f[439] && f[521] && f[304] && !f[382]; // c8t108i10
	assign leaf[175] = f[439] && f[521] && f[304] && f[382]; // c8t108i10
	assign leaf[176] = !f[438] && !f[434] && !f[378] && !f[410]; // c8t118i11
	assign leaf[177] = !f[438] && !f[434] && !f[378] && f[410]; // c8t118i11
	assign leaf[178] = !f[438] && !f[434] && f[378] && !f[153]; // c8t118i11
	assign leaf[179] = !f[438] && !f[434] && f[378] && f[153]; // c8t118i11
	assign leaf[180] = !f[438] && f[434] && !f[687] && !f[292]; // c8t118i11
	assign leaf[181] = !f[438] && f[434] && !f[687] && f[292]; // c8t118i11
	assign leaf[182] = !f[438] && f[434] && f[687] && !f[544]; // c8t118i11
	assign leaf[183] = !f[438] && f[434] && f[687] && f[544]; // c8t118i11
	assign leaf[184] = f[438] && !f[520] && !f[330] && !f[153]; // c8t118i11
	assign leaf[185] = f[438] && !f[520] && !f[330] && f[153]; // c8t118i11
	assign leaf[186] = f[438] && !f[520] && f[330] && !f[300]; // c8t118i11
	assign leaf[187] = f[438] && !f[520] && f[330] && f[300]; // c8t118i11
	assign leaf[188] = f[438] && f[520] && !f[302] && !f[331]; // c8t118i11
	assign leaf[189] = f[438] && f[520] && !f[302] && f[331]; // c8t118i11
	assign leaf[190] = f[438] && f[520] && f[302] && !f[427]; // c8t118i11
	assign leaf[191] = f[438] && f[520] && f[302] && f[427]; // c8t118i11
	assign leaf[192] = !f[274] && !f[660] && !f[597] && !f[567]; // c8t128i12
	assign leaf[193] = !f[274] && !f[660] && !f[597] && f[567]; // c8t128i12
	assign leaf[194] = !f[274] && !f[660] && f[597] && !f[572]; // c8t128i12
	assign leaf[195] = !f[274] && !f[660] && f[597] && f[572]; // c8t128i12
	assign leaf[196] = !f[274] && f[660] && !f[544] && !f[542]; // c8t128i12
	assign leaf[197] = !f[274] && f[660] && !f[544] && f[542]; // c8t128i12
	assign leaf[198] = !f[274] && f[660] && f[544] && !f[513]; // c8t128i12
	assign leaf[199] = !f[274] && f[660] && f[544] && f[513]; // c8t128i12
	assign leaf[200] = f[274] && !f[426] && !f[271] && !f[380]; // c8t128i12
	assign leaf[201] = f[274] && !f[426] && !f[271] && f[380]; // c8t128i12
	assign leaf[202] = f[274] && !f[426] && f[271] && !f[486]; // c8t128i12
	assign leaf[203] = f[274] && !f[426] && f[271] && f[486]; // c8t128i12
	assign leaf[204] = f[274] && f[426] && !f[520] && !f[409]; // c8t128i12
	assign leaf[205] = f[274] && f[426] && !f[520] && f[409]; // c8t128i12
	assign leaf[206] = f[274] && f[426] && f[520] && !f[634]; // c8t128i12
	assign leaf[207] = f[274] && f[426] && f[520] && f[634]; // c8t128i12
	assign leaf[208] = !f[440] && !f[288] && !f[541] && !f[511]; // c8t138i13
	assign leaf[209] = !f[440] && !f[288] && !f[541] && f[511]; // c8t138i13
	assign leaf[210] = !f[440] && !f[288] && f[541] && !f[571]; // c8t138i13
	assign leaf[211] = !f[440] && !f[288] && f[541] && f[571]; // c8t138i13
	assign leaf[212] = !f[440] && f[288] && !f[374] && !f[348]; // c8t138i13
	assign leaf[213] = !f[440] && f[288] && !f[374] && f[348]; // c8t138i13
	assign leaf[214] = !f[440] && f[288] && f[374] && !f[517]; // c8t138i13
	assign leaf[215] = !f[440] && f[288] && f[374] && f[517]; // c8t138i13
	assign leaf[216] = f[440] && !f[582] && !f[304] && !f[494]; // c8t138i13
	assign leaf[217] = f[440] && !f[582] && !f[304] && f[494]; // c8t138i13
	assign leaf[218] = f[440] && !f[582] && f[304] && !f[371]; // c8t138i13
	assign leaf[219] = f[440] && !f[582] && f[304] && f[371]; // c8t138i13
	assign leaf[220] = f[440] && f[582] && !f[525] && !f[349]; // c8t138i13
	assign leaf[221] = f[440] && f[582] && !f[525] && f[349]; // c8t138i13
	assign leaf[222] = f[440] && f[582] && f[525] && !f[460]; // c8t138i13
	assign leaf[223] = f[440] && f[582] && f[525] && f[460]; // c8t138i13
	assign leaf[224] = !f[466] && !f[185] && !f[157] && !f[627]; // c8t148i14
	assign leaf[225] = !f[466] && !f[185] && !f[157] && f[627]; // c8t148i14
	assign leaf[226] = !f[466] && !f[185] && f[157] && !f[580]; // c8t148i14
	assign leaf[227] = !f[466] && !f[185] && f[157] && f[580]; // c8t148i14
	assign leaf[228] = !f[466] && f[185] && !f[268] && !f[322]; // c8t148i14
	assign leaf[229] = !f[466] && f[185] && !f[268] && f[322]; // c8t148i14
	assign leaf[230] = !f[466] && f[185] && f[268] && !f[659]; // c8t148i14
	assign leaf[231] = !f[466] && f[185] && f[268] && f[659]; // c8t148i14
	assign leaf[232] = f[466] && !f[520] && !f[350] && !f[233]; // c8t148i14
	assign leaf[233] = f[466] && !f[520] && !f[350] && f[233]; // c8t148i14
	assign leaf[234] = f[466] && !f[520] && f[350] && !f[440]; // c8t148i14
	assign leaf[235] = f[466] && !f[520] && f[350] && f[440]; // c8t148i14
	assign leaf[236] = f[466] && f[520] && !f[180] && !f[620]; // c8t148i14
	assign leaf[237] = f[466] && f[520] && !f[180] && f[620]; // c8t148i14
	assign leaf[238] = f[466] && f[520] && f[180] && !f[275]; // c8t148i14
	assign leaf[239] = f[466] && f[520] && f[180] && f[275]; // c8t148i14
	assign leaf[240] = !f[467] && !f[658] && !f[513] && !f[663]; // c8t158i15
	assign leaf[241] = !f[467] && !f[658] && !f[513] && f[663]; // c8t158i15
	assign leaf[242] = !f[467] && !f[658] && f[513] && !f[628]; // c8t158i15
	assign leaf[243] = !f[467] && !f[658] && f[513] && f[628]; // c8t158i15
	assign leaf[244] = !f[467] && f[658] && !f[602] && !f[572]; // c8t158i15
	assign leaf[245] = !f[467] && f[658] && !f[602] && f[572]; // c8t158i15
	assign leaf[246] = !f[467] && f[658] && f[602] && !f[267]; // c8t158i15
	assign leaf[247] = !f[467] && f[658] && f[602] && f[267]; // c8t158i15
	assign leaf[248] = f[467] && !f[521] && !f[638] && !f[261]; // c8t158i15
	assign leaf[249] = f[467] && !f[521] && !f[638] && f[261]; // c8t158i15
	assign leaf[250] = f[467] && !f[521] && f[638] && !f[551]; // c8t158i15
	assign leaf[251] = f[467] && !f[521] && f[638] && f[551]; // c8t158i15
	assign leaf[252] = f[467] && f[521] && !f[351] && !f[637]; // c8t158i15
	assign leaf[253] = f[467] && f[521] && !f[351] && f[637]; // c8t158i15
	assign leaf[254] = f[467] && f[521] && f[351] && !f[274]; // c8t158i15
	assign leaf[255] = f[467] && f[521] && f[351] && f[274]; // c8t158i15
	assign leaf[256] = !f[434] && !f[520] && !f[549] && !f[457]; // c8t168i16
	assign leaf[257] = !f[434] && !f[520] && !f[549] && f[457]; // c8t168i16
	assign leaf[258] = !f[434] && !f[520] && f[549] && !f[407]; // c8t168i16
	assign leaf[259] = !f[434] && !f[520] && f[549] && f[407]; // c8t168i16
	assign leaf[260] = !f[434] && f[520] && !f[378] && !f[304]; // c8t168i16
	assign leaf[261] = !f[434] && f[520] && !f[378] && f[304]; // c8t168i16
	assign leaf[262] = !f[434] && f[520] && f[378] && !f[346]; // c8t168i16
	assign leaf[263] = !f[434] && f[520] && f[378] && f[346]; // c8t168i16
	assign leaf[264] = f[434] && !f[437] && !f[124] && !f[496]; // c8t168i16
	assign leaf[265] = f[434] && !f[437] && !f[124] && f[496]; // c8t168i16
	assign leaf[266] = f[434] && !f[437] && f[124] && !f[465]; // c8t168i16
	assign leaf[267] = f[434] && !f[437] && f[124] && f[465]; // c8t168i16
	assign leaf[268] = f[434] && f[437] && !f[634] && !f[541]; // c8t168i16
	assign leaf[269] = f[434] && f[437] && !f[634] && f[541]; // c8t168i16
	assign leaf[270] = f[434] && f[437] && f[634] && !f[315]; // c8t168i16
	assign leaf[271] = f[434] && f[437] && f[634] && f[315]; // c8t168i16
	assign leaf[272] = !f[440] && !f[357] && !f[410] && !f[289]; // c8t178i17
	assign leaf[273] = !f[440] && !f[357] && !f[410] && f[289]; // c8t178i17
	assign leaf[274] = !f[440] && !f[357] && f[410] && !f[465]; // c8t178i17
	assign leaf[275] = !f[440] && !f[357] && f[410] && f[465]; // c8t178i17
	assign leaf[276] = !f[440] && f[357] && !f[327] && !f[469]; // c8t178i17
	assign leaf[277] = !f[440] && f[357] && !f[327] && f[469]; // c8t178i17
	assign leaf[278] = !f[440] && f[357] && f[327] && !f[185]; // c8t178i17
	assign leaf[279] = !f[440] && f[357] && f[327] && f[185]; // c8t178i17
	assign leaf[280] = f[440] && !f[522] && !f[180] && !f[360]; // c8t178i17
	assign leaf[281] = f[440] && !f[522] && !f[180] && f[360]; // c8t178i17
	assign leaf[282] = f[440] && !f[522] && f[180] && !f[210]; // c8t178i17
	assign leaf[283] = f[440] && !f[522] && f[180] && f[210]; // c8t178i17
	assign leaf[284] = f[440] && f[522] && !f[303] && !f[611]; // c8t178i17
	assign leaf[285] = f[440] && f[522] && !f[303] && f[611]; // c8t178i17
	assign leaf[286] = f[440] && f[522] && f[303] && !f[399]; // c8t178i17
	assign leaf[287] = f[440] && f[522] && f[303] && f[399]; // c8t178i17
	assign leaf[288] = !f[434] && !f[520] && !f[457] && !f[459]; // c8t188i18
	assign leaf[289] = !f[434] && !f[520] && !f[457] && f[459]; // c8t188i18
	assign leaf[290] = !f[434] && !f[520] && f[457] && !f[380]; // c8t188i18
	assign leaf[291] = !f[434] && !f[520] && f[457] && f[380]; // c8t188i18
	assign leaf[292] = !f[434] && f[520] && !f[347] && !f[459]; // c8t188i18
	assign leaf[293] = !f[434] && f[520] && !f[347] && f[459]; // c8t188i18
	assign leaf[294] = !f[434] && f[520] && f[347] && !f[378]; // c8t188i18
	assign leaf[295] = !f[434] && f[520] && f[347] && f[378]; // c8t188i18
	assign leaf[296] = f[434] && !f[428] && !f[316] && !f[291]; // c8t188i18
	assign leaf[297] = f[434] && !f[428] && !f[316] && f[291]; // c8t188i18
	assign leaf[298] = f[434] && !f[428] && f[316] && !f[374]; // c8t188i18
	assign leaf[299] = f[434] && !f[428] && f[316] && f[374]; // c8t188i18
	assign leaf[300] = f[434] && f[428] && !f[662] && !f[595]; // c8t188i18
	assign leaf[301] = f[434] && f[428] && !f[662] && f[595]; // c8t188i18
	assign leaf[302] = f[434] && f[428] && f[662] && !f[573]; // c8t188i18
	assign leaf[303] = f[434] && f[428] && f[662] && f[573]; // c8t188i18
	assign leaf[304] = !f[302] && !f[332] && !f[349] && !f[375]; // c8t198i19
	assign leaf[305] = !f[302] && !f[332] && !f[349] && f[375]; // c8t198i19
	assign leaf[306] = !f[302] && !f[332] && f[349] && !f[375]; // c8t198i19
	assign leaf[307] = !f[302] && !f[332] && f[349] && f[375]; // c8t198i19
	assign leaf[308] = !f[302] && f[332] && !f[385]; // c8t198i19
	assign leaf[309] = !f[302] && f[332] && f[385] && !f[653]; // c8t198i19
	assign leaf[310] = !f[302] && f[332] && f[385] && f[653]; // c8t198i19
	assign leaf[311] = f[302] && !f[272] && !f[399] && !f[601]; // c8t198i19
	assign leaf[312] = f[302] && !f[272] && !f[399] && f[601]; // c8t198i19
	assign leaf[313] = f[302] && !f[272] && f[399] && !f[687]; // c8t198i19
	assign leaf[314] = f[302] && !f[272] && f[399] && f[687]; // c8t198i19
	assign leaf[315] = f[302] && f[272] && !f[458] && !f[296]; // c8t198i19
	assign leaf[316] = f[302] && f[272] && !f[458] && f[296]; // c8t198i19
	assign leaf[317] = f[302] && f[272] && f[458] && !f[352]; // c8t198i19
	assign leaf[318] = f[302] && f[272] && f[458] && f[352]; // c8t198i19
	assign leaf[319] = !f[441] && !f[314] && !f[401] && !f[318]; // c8t208i20
	assign leaf[320] = !f[441] && !f[314] && !f[401] && f[318]; // c8t208i20
	assign leaf[321] = !f[441] && !f[314] && f[401] && !f[437]; // c8t208i20
	assign leaf[322] = !f[441] && !f[314] && f[401] && f[437]; // c8t208i20
	assign leaf[323] = !f[441] && f[314] && !f[402] && !f[375]; // c8t208i20
	assign leaf[324] = !f[441] && f[314] && !f[402] && f[375]; // c8t208i20
	assign leaf[325] = !f[441] && f[314] && f[402] && !f[517]; // c8t208i20
	assign leaf[326] = !f[441] && f[314] && f[402] && f[517]; // c8t208i20
	assign leaf[327] = f[441] && !f[523] && !f[595] && !f[608]; // c8t208i20
	assign leaf[328] = f[441] && !f[523] && !f[595] && f[608]; // c8t208i20
	assign leaf[329] = f[441] && !f[523] && f[595] && !f[403]; // c8t208i20
	assign leaf[330] = f[441] && !f[523] && f[595] && f[403]; // c8t208i20
	assign leaf[331] = f[441] && f[523] && !f[593] && !f[691]; // c8t208i20
	assign leaf[332] = f[441] && f[523] && !f[593] && f[691]; // c8t208i20
	assign leaf[333] = f[441] && f[523] && f[593] && !f[330]; // c8t208i20
	assign leaf[334] = f[441] && f[523] && f[593] && f[330]; // c8t208i20
	assign leaf[335] = !f[153] && !f[186] && !f[158] && !f[542]; // c8t218i21
	assign leaf[336] = !f[153] && !f[186] && !f[158] && f[542]; // c8t218i21
	assign leaf[337] = !f[153] && !f[186] && f[158] && !f[326]; // c8t218i21
	assign leaf[338] = !f[153] && !f[186] && f[158] && f[326]; // c8t218i21
	assign leaf[339] = !f[153] && f[186] && !f[241] && !f[322]; // c8t218i21
	assign leaf[340] = !f[153] && f[186] && !f[241] && f[322]; // c8t218i21
	assign leaf[341] = !f[153] && f[186] && f[241] && !f[659]; // c8t218i21
	assign leaf[342] = !f[153] && f[186] && f[241] && f[659]; // c8t218i21
	assign leaf[343] = f[153] && !f[210] && !f[350] && !f[376]; // c8t218i21
	assign leaf[344] = f[153] && !f[210] && !f[350] && f[376]; // c8t218i21
	assign leaf[345] = f[153] && !f[210] && f[350] && !f[293]; // c8t218i21
	assign leaf[346] = f[153] && !f[210] && f[350] && f[293]; // c8t218i21
	assign leaf[347] = f[153] && f[210] && !f[289] && !f[343]; // c8t218i21
	assign leaf[348] = f[153] && f[210] && !f[289] && f[343]; // c8t218i21
	assign leaf[349] = f[153] && f[210] && f[289] && !f[264]; // c8t218i21
	assign leaf[350] = f[153] && f[210] && f[289] && f[264]; // c8t218i21
	assign leaf[351] = !f[688] && !f[219] && !f[631] && !f[596]; // c8t228i22
	assign leaf[352] = !f[688] && !f[219] && !f[631] && f[596]; // c8t228i22
	assign leaf[353] = !f[688] && !f[219] && f[631] && !f[516]; // c8t228i22
	assign leaf[354] = !f[688] && !f[219] && f[631] && f[516]; // c8t228i22
	assign leaf[355] = !f[688] && f[219] && !f[400] && !f[508]; // c8t228i22
	assign leaf[356] = !f[688] && f[219] && !f[400] && f[508]; // c8t228i22
	assign leaf[357] = !f[688] && f[219] && f[400] && !f[347]; // c8t228i22
	assign leaf[358] = !f[688] && f[219] && f[400] && f[347]; // c8t228i22
	assign leaf[359] = f[688] && !f[573] && !f[571] && !f[569]; // c8t228i22
	assign leaf[360] = f[688] && !f[573] && !f[571] && f[569]; // c8t228i22
	assign leaf[361] = f[688] && !f[573] && f[571] && !f[630]; // c8t228i22
	assign leaf[362] = f[688] && !f[573] && f[571] && f[630]; // c8t228i22
	assign leaf[363] = f[688] && f[573] && !f[513] && !f[717]; // c8t228i22
	assign leaf[364] = f[688] && f[573] && !f[513] && f[717]; // c8t228i22
	assign leaf[365] = f[688] && f[573] && f[513] && !f[214]; // c8t228i22
	assign leaf[366] = f[688] && f[573] && f[513] && f[214]; // c8t228i22
	assign leaf[367] = !f[301] && !f[330] && !f[271] && !f[300]; // c8t238i23
	assign leaf[368] = !f[301] && !f[330] && !f[271] && f[300]; // c8t238i23
	assign leaf[369] = !f[301] && !f[330] && f[271] && !f[242]; // c8t238i23
	assign leaf[370] = !f[301] && !f[330] && f[271] && f[242]; // c8t238i23
	assign leaf[371] = !f[301] && f[330] && !f[524] && !f[439]; // c8t238i23
	assign leaf[372] = !f[301] && f[330] && !f[524] && f[439]; // c8t238i23
	assign leaf[373] = !f[301] && f[330] && f[524]; // c8t238i23
	assign leaf[374] = f[301] && !f[298] && !f[322] && !f[399]; // c8t238i23
	assign leaf[375] = f[301] && !f[298] && !f[322] && f[399]; // c8t238i23
	assign leaf[376] = f[301] && !f[298] && f[322] && !f[536]; // c8t238i23
	assign leaf[377] = f[301] && !f[298] && f[322] && f[536]; // c8t238i23
	assign leaf[378] = f[301] && f[298] && !f[458] && !f[459]; // c8t238i23
	assign leaf[379] = f[301] && f[298] && !f[458] && f[459]; // c8t238i23
	assign leaf[380] = f[301] && f[298] && f[458] && !f[243]; // c8t238i23
	assign leaf[381] = f[301] && f[298] && f[458] && f[243]; // c8t238i23
	assign leaf[382] = !f[322] && !f[489] && !f[487] && !f[484]; // c8t248i24
	assign leaf[383] = !f[322] && !f[489] && !f[487] && f[484]; // c8t248i24
	assign leaf[384] = !f[322] && !f[489] && f[487] && !f[457]; // c8t248i24
	assign leaf[385] = !f[322] && !f[489] && f[487] && f[457]; // c8t248i24
	assign leaf[386] = !f[322] && f[489] && !f[376] && !f[402]; // c8t248i24
	assign leaf[387] = !f[322] && f[489] && !f[376] && f[402]; // c8t248i24
	assign leaf[388] = !f[322] && f[489] && f[376] && !f[430]; // c8t248i24
	assign leaf[389] = !f[322] && f[489] && f[376] && f[430]; // c8t248i24
	assign leaf[390] = f[322] && !f[239] && !f[155] && !f[602]; // c8t248i24
	assign leaf[391] = f[322] && !f[239] && !f[155] && f[602]; // c8t248i24
	assign leaf[392] = f[322] && !f[239] && f[155] && !f[293]; // c8t248i24
	assign leaf[393] = f[322] && !f[239] && f[155] && f[293]; // c8t248i24
	assign leaf[394] = f[322] && f[239] && !f[296] && !f[348]; // c8t248i24
	assign leaf[395] = f[322] && f[239] && !f[296] && f[348]; // c8t248i24
	assign leaf[396] = f[322] && f[239] && f[296] && !f[662]; // c8t248i24
	assign leaf[397] = f[322] && f[239] && f[296] && f[662]; // c8t248i24
	assign leaf[398] = !f[287] && !f[468] && !f[357] && !f[410]; // c8t258i25
	assign leaf[399] = !f[287] && !f[468] && !f[357] && f[410]; // c8t258i25
	assign leaf[400] = !f[287] && !f[468] && f[357] && !f[327]; // c8t258i25
	assign leaf[401] = !f[287] && !f[468] && f[357] && f[327]; // c8t258i25
	assign leaf[402] = !f[287] && f[468] && !f[322] && !f[354]; // c8t258i25
	assign leaf[403] = !f[287] && f[468] && !f[322] && f[354]; // c8t258i25
	assign leaf[404] = !f[287] && f[468] && f[322] && !f[262]; // c8t258i25
	assign leaf[405] = !f[287] && f[468] && f[322] && f[262]; // c8t258i25
	assign leaf[406] = f[287] && !f[517] && !f[346] && !f[401]; // c8t258i25
	assign leaf[407] = f[287] && !f[517] && !f[346] && f[401]; // c8t258i25
	assign leaf[408] = f[287] && !f[517] && f[346] && !f[371]; // c8t258i25
	assign leaf[409] = f[287] && !f[517] && f[346] && f[371]; // c8t258i25
	assign leaf[410] = f[287] && f[517] && !f[514] && !f[682]; // c8t258i25
	assign leaf[411] = f[287] && f[517] && !f[514] && f[682]; // c8t258i25
	assign leaf[412] = f[287] && f[517] && f[514] && !f[343]; // c8t258i25
	assign leaf[413] = f[287] && f[517] && f[514] && f[343]; // c8t258i25
	assign leaf[414] = !f[469] && !f[287] && !f[274] && !f[330]; // c8t268i26
	assign leaf[415] = !f[469] && !f[287] && !f[274] && f[330]; // c8t268i26
	assign leaf[416] = !f[469] && !f[287] && f[274] && !f[677]; // c8t268i26
	assign leaf[417] = !f[469] && !f[287] && f[274] && f[677]; // c8t268i26
	assign leaf[418] = !f[469] && f[287] && !f[374] && !f[400]; // c8t268i26
	assign leaf[419] = !f[469] && f[287] && !f[374] && f[400]; // c8t268i26
	assign leaf[420] = !f[469] && f[287] && f[374] && !f[438]; // c8t268i26
	assign leaf[421] = !f[469] && f[287] && f[374] && f[438]; // c8t268i26
	assign leaf[422] = f[469] && !f[523] && !f[206] && !f[570]; // c8t268i26
	assign leaf[423] = f[469] && !f[523] && !f[206] && f[570]; // c8t268i26
	assign leaf[424] = f[469] && !f[523] && f[206] && !f[401]; // c8t268i26
	assign leaf[425] = f[469] && !f[523] && f[206] && f[401]; // c8t268i26
	assign leaf[426] = f[469] && f[523] && !f[569] && !f[161]; // c8t268i26
	assign leaf[427] = f[469] && f[523] && !f[569] && f[161]; // c8t268i26
	assign leaf[428] = f[469] && f[523] && f[569] && !f[414]; // c8t268i26
	assign leaf[429] = f[469] && f[523] && f[569] && f[414]; // c8t268i26
	assign leaf[430] = !f[441] && !f[314] && !f[437] && !f[406]; // c8t278i27
	assign leaf[431] = !f[441] && !f[314] && !f[437] && f[406]; // c8t278i27
	assign leaf[432] = !f[441] && !f[314] && f[437] && !f[152]; // c8t278i27
	assign leaf[433] = !f[441] && !f[314] && f[437] && f[152]; // c8t278i27
	assign leaf[434] = !f[441] && f[314] && !f[353] && !f[296]; // c8t278i27
	assign leaf[435] = !f[441] && f[314] && !f[353] && f[296]; // c8t278i27
	assign leaf[436] = !f[441] && f[314] && f[353] && !f[431]; // c8t278i27
	assign leaf[437] = !f[441] && f[314] && f[353] && f[431]; // c8t278i27
	assign leaf[438] = f[441] && !f[332] && !f[555] && !f[593]; // c8t278i27
	assign leaf[439] = f[441] && !f[332] && !f[555] && f[593]; // c8t278i27
	assign leaf[440] = f[441] && !f[332] && f[555] && !f[300]; // c8t278i27
	assign leaf[441] = f[441] && !f[332] && f[555] && f[300]; // c8t278i27
	assign leaf[442] = f[441] && f[332] && !f[549] && !f[187]; // c8t278i27
	assign leaf[443] = f[441] && f[332] && !f[549] && f[187]; // c8t278i27
	assign leaf[444] = f[441] && f[332] && f[549]; // c8t278i27
	assign leaf[445] = !f[322] && !f[489] && !f[663] && !f[301]; // c8t288i28
	assign leaf[446] = !f[322] && !f[489] && !f[663] && f[301]; // c8t288i28
	assign leaf[447] = !f[322] && !f[489] && f[663] && !f[546]; // c8t288i28
	assign leaf[448] = !f[322] && !f[489] && f[663] && f[546]; // c8t288i28
	assign leaf[449] = !f[322] && f[489] && !f[485] && !f[659]; // c8t288i28
	assign leaf[450] = !f[322] && f[489] && !f[485] && f[659]; // c8t288i28
	assign leaf[451] = !f[322] && f[489] && f[485] && !f[493]; // c8t288i28
	assign leaf[452] = !f[322] && f[489] && f[485] && f[493]; // c8t288i28
	assign leaf[453] = f[322] && !f[546] && !f[264] && !f[290]; // c8t288i28
	assign leaf[454] = f[322] && !f[546] && !f[264] && f[290]; // c8t288i28
	assign leaf[455] = f[322] && !f[546] && f[264] && !f[238]; // c8t288i28
	assign leaf[456] = f[322] && !f[546] && f[264] && f[238]; // c8t288i28
	assign leaf[457] = f[322] && f[546] && !f[348] && !f[296]; // c8t288i28
	assign leaf[458] = f[322] && f[546] && !f[348] && f[296]; // c8t288i28
	assign leaf[459] = f[322] && f[546] && f[348] && !f[233]; // c8t288i28
	assign leaf[460] = f[322] && f[546] && f[348] && f[233]; // c8t288i28
	assign leaf[461] = !f[261] && !f[374] && !f[292] && !f[266]; // c8t298i29
	assign leaf[462] = !f[261] && !f[374] && !f[292] && f[266]; // c8t298i29
	assign leaf[463] = !f[261] && !f[374] && f[292] && !f[238]; // c8t298i29
	assign leaf[464] = !f[261] && !f[374] && f[292] && f[238]; // c8t298i29
	assign leaf[465] = !f[261] && f[374] && !f[286] && !f[320]; // c8t298i29
	assign leaf[466] = !f[261] && f[374] && !f[286] && f[320]; // c8t298i29
	assign leaf[467] = !f[261] && f[374] && f[286] && !f[398]; // c8t298i29
	assign leaf[468] = !f[261] && f[374] && f[286] && f[398]; // c8t298i29
	assign leaf[469] = f[261] && !f[348] && !f[374] && !f[401]; // c8t298i29
	assign leaf[470] = f[261] && !f[348] && !f[374] && f[401]; // c8t298i29
	assign leaf[471] = f[261] && !f[348] && f[374] && !f[489]; // c8t298i29
	assign leaf[472] = f[261] && !f[348] && f[374] && f[489]; // c8t298i29
	assign leaf[473] = f[261] && f[348] && !f[372] && !f[235]; // c8t298i29
	assign leaf[474] = f[261] && f[348] && !f[372] && f[235]; // c8t298i29
	assign leaf[475] = f[261] && f[348] && f[372] && !f[434]; // c8t298i29
	assign leaf[476] = f[261] && f[348] && f[372] && f[434]; // c8t298i29
	assign leaf[477] = !f[219] && !f[467] && !f[315] && !f[202]; // c8t308i30
	assign leaf[478] = !f[219] && !f[467] && !f[315] && f[202]; // c8t308i30
	assign leaf[479] = !f[219] && !f[467] && f[315] && !f[290]; // c8t308i30
	assign leaf[480] = !f[219] && !f[467] && f[315] && f[290]; // c8t308i30
	assign leaf[481] = !f[219] && f[467] && !f[521] && !f[638]; // c8t308i30
	assign leaf[482] = !f[219] && f[467] && !f[521] && f[638]; // c8t308i30
	assign leaf[483] = !f[219] && f[467] && f[521] && !f[637]; // c8t308i30
	assign leaf[484] = !f[219] && f[467] && f[521] && f[637]; // c8t308i30
	assign leaf[485] = f[219] && !f[458] && !f[655] && !f[685]; // c8t308i30
	assign leaf[486] = f[219] && !f[458] && !f[655] && f[685]; // c8t308i30
	assign leaf[487] = f[219] && !f[458] && f[655] && !f[346]; // c8t308i30
	assign leaf[488] = f[219] && !f[458] && f[655] && f[346]; // c8t308i30
	assign leaf[489] = f[219] && f[458] && !f[460] && !f[247]; // c8t308i30
	assign leaf[490] = f[219] && f[458] && !f[460] && f[247]; // c8t308i30
	assign leaf[491] = f[219] && f[458] && f[460] && !f[428]; // c8t308i30
	assign leaf[492] = f[219] && f[458] && f[460] && f[428]; // c8t308i30
	assign leaf[493] = !f[439] && !f[525] && !f[542] && !f[512]; // c8t318i31
	assign leaf[494] = !f[439] && !f[525] && !f[542] && f[512]; // c8t318i31
	assign leaf[495] = !f[439] && !f[525] && f[542] && !f[544]; // c8t318i31
	assign leaf[496] = !f[439] && !f[525] && f[542] && f[544]; // c8t318i31
	assign leaf[497] = !f[439] && f[525] && !f[637] && !f[383]; // c8t318i31
	assign leaf[498] = !f[439] && f[525] && !f[637] && f[383]; // c8t318i31
	assign leaf[499] = !f[439] && f[525] && f[637] && !f[377]; // c8t318i31
	assign leaf[500] = !f[439] && f[525] && f[637] && f[377]; // c8t318i31
	assign leaf[501] = f[439] && !f[521] && !f[271] && !f[217]; // c8t318i31
	assign leaf[502] = f[439] && !f[521] && !f[271] && f[217]; // c8t318i31
	assign leaf[503] = f[439] && !f[521] && f[271] && !f[298]; // c8t318i31
	assign leaf[504] = f[439] && !f[521] && f[271] && f[298]; // c8t318i31
	assign leaf[505] = f[439] && f[521] && !f[594] && !f[153]; // c8t318i31
	assign leaf[506] = f[439] && f[521] && !f[594] && f[153]; // c8t318i31
	assign leaf[507] = f[439] && f[521] && f[594] && !f[457]; // c8t318i31
	assign leaf[508] = f[439] && f[521] && f[594] && f[457]; // c8t318i31
	assign leaf[509] = !f[441] && !f[341] && !f[357] && !f[410]; // c8t328i32
	assign leaf[510] = !f[441] && !f[341] && !f[357] && f[410]; // c8t328i32
	assign leaf[511] = !f[441] && !f[341] && f[357] && !f[328]; // c8t328i32
	assign leaf[512] = !f[441] && !f[341] && f[357] && f[328]; // c8t328i32
	assign leaf[513] = !f[441] && f[341] && !f[315] && !f[430]; // c8t328i32
	assign leaf[514] = !f[441] && f[341] && !f[315] && f[430]; // c8t328i32
	assign leaf[515] = !f[441] && f[341] && f[315] && !f[435]; // c8t328i32
	assign leaf[516] = !f[441] && f[341] && f[315] && f[435]; // c8t328i32
	assign leaf[517] = f[441] && !f[595] && !f[523] && !f[633]; // c8t328i32
	assign leaf[518] = f[441] && !f[595] && !f[523] && f[633]; // c8t328i32
	assign leaf[519] = f[441] && !f[595] && f[523] && !f[691]; // c8t328i32
	assign leaf[520] = f[441] && !f[595] && f[523] && f[691]; // c8t328i32
	assign leaf[521] = f[441] && f[595] && !f[496] && !f[510]; // c8t328i32
	assign leaf[522] = f[441] && f[595] && !f[496] && f[510]; // c8t328i32
	assign leaf[523] = f[441] && f[595] && f[496] && !f[456]; // c8t328i32
	assign leaf[524] = f[441] && f[595] && f[496] && f[456]; // c8t328i32
	assign leaf[525] = !f[440] && !f[315] && !f[290] && !f[292]; // c8t338i33
	assign leaf[526] = !f[440] && !f[315] && !f[290] && f[292]; // c8t338i33
	assign leaf[527] = !f[440] && !f[315] && f[290] && !f[264]; // c8t338i33
	assign leaf[528] = !f[440] && !f[315] && f[290] && f[264]; // c8t338i33
	assign leaf[529] = !f[440] && f[315] && !f[489] && !f[288]; // c8t338i33
	assign leaf[530] = !f[440] && f[315] && !f[489] && f[288]; // c8t338i33
	assign leaf[531] = !f[440] && f[315] && f[489] && !f[634]; // c8t338i33
	assign leaf[532] = !f[440] && f[315] && f[489] && f[634]; // c8t338i33
	assign leaf[533] = f[440] && !f[576] && !f[567] && !f[514]; // c8t338i33
	assign leaf[534] = f[440] && !f[576] && !f[567] && f[514]; // c8t338i33
	assign leaf[535] = f[440] && !f[576] && f[567] && !f[681]; // c8t338i33
	assign leaf[536] = f[440] && !f[576] && f[567] && f[681]; // c8t338i33
	assign leaf[537] = f[440] && f[576] && !f[637] && !f[634]; // c8t338i33
	assign leaf[538] = f[440] && f[576] && !f[637] && f[634]; // c8t338i33
	assign leaf[539] = f[440] && f[576] && f[637] && !f[657]; // c8t338i33
	assign leaf[540] = f[440] && f[576] && f[637] && f[657]; // c8t338i33
	assign leaf[541] = !f[248] && !f[350] && !f[517] && !f[514]; // c8t348i34
	assign leaf[542] = !f[248] && !f[350] && !f[517] && f[514]; // c8t348i34
	assign leaf[543] = !f[248] && !f[350] && f[517] && !f[456]; // c8t348i34
	assign leaf[544] = !f[248] && !f[350] && f[517] && f[456]; // c8t348i34
	assign leaf[545] = !f[248] && f[350] && !f[517] && !f[293]; // c8t348i34
	assign leaf[546] = !f[248] && f[350] && !f[517] && f[293]; // c8t348i34
	assign leaf[547] = !f[248] && f[350] && f[517] && !f[632]; // c8t348i34
	assign leaf[548] = !f[248] && f[350] && f[517] && f[632]; // c8t348i34
	assign leaf[549] = f[248] && !f[186] && !f[401] && !f[485]; // c8t348i34
	assign leaf[550] = f[248] && !f[186] && !f[401] && f[485]; // c8t348i34
	assign leaf[551] = f[248] && !f[186] && f[401] && !f[432]; // c8t348i34
	assign leaf[552] = f[248] && !f[186] && f[401] && f[432]; // c8t348i34
	assign leaf[553] = f[248] && f[186] && !f[577] && !f[181]; // c8t348i34
	assign leaf[554] = f[248] && f[186] && !f[577] && f[181]; // c8t348i34
	assign leaf[555] = f[248] && f[186] && f[577] && !f[328]; // c8t348i34
	assign leaf[556] = f[248] && f[186] && f[577] && f[328]; // c8t348i34
	assign leaf[557] = !f[248] && !f[156] && !f[542] && !f[544]; // c8t358i35
	assign leaf[558] = !f[248] && !f[156] && !f[542] && f[544]; // c8t358i35
	assign leaf[559] = !f[248] && !f[156] && f[542] && !f[455]; // c8t358i35
	assign leaf[560] = !f[248] && !f[156] && f[542] && f[455]; // c8t358i35
	assign leaf[561] = !f[248] && f[156] && !f[212] && !f[266]; // c8t358i35
	assign leaf[562] = !f[248] && f[156] && !f[212] && f[266]; // c8t358i35
	assign leaf[563] = !f[248] && f[156] && f[212] && !f[576]; // c8t358i35
	assign leaf[564] = !f[248] && f[156] && f[212] && f[576]; // c8t358i35
	assign leaf[565] = f[248] && !f[347] && !f[322] && !f[575]; // c8t358i35
	assign leaf[566] = f[248] && !f[347] && !f[322] && f[575]; // c8t358i35
	assign leaf[567] = f[248] && !f[347] && f[322] && !f[352]; // c8t358i35
	assign leaf[568] = f[248] && !f[347] && f[322] && f[352]; // c8t358i35
	assign leaf[569] = f[248] && f[347] && !f[383] && !f[374]; // c8t358i35
	assign leaf[570] = f[248] && f[347] && !f[383] && f[374]; // c8t358i35
	assign leaf[571] = f[248] && f[347] && f[383] && !f[371]; // c8t358i35
	assign leaf[572] = f[248] && f[347] && f[383] && f[371]; // c8t358i35
	assign leaf[573] = !f[340] && !f[399] && !f[317] && !f[291]; // c8t368i36
	assign leaf[574] = !f[340] && !f[399] && !f[317] && f[291]; // c8t368i36
	assign leaf[575] = !f[340] && !f[399] && f[317] && !f[403]; // c8t368i36
	assign leaf[576] = !f[340] && !f[399] && f[317] && f[403]; // c8t368i36
	assign leaf[577] = !f[340] && f[399] && !f[493] && !f[510]; // c8t368i36
	assign leaf[578] = !f[340] && f[399] && !f[493] && f[510]; // c8t368i36
	assign leaf[579] = !f[340] && f[399] && f[493] && !f[346]; // c8t368i36
	assign leaf[580] = !f[340] && f[399] && f[493] && f[346]; // c8t368i36
	assign leaf[581] = f[340] && !f[464]; // c8t368i36
	assign leaf[582] = f[340] && f[464] && !f[152] && !f[546]; // c8t368i36
	assign leaf[583] = f[340] && f[464] && !f[152] && f[546]; // c8t368i36
	assign leaf[584] = f[340] && f[464] && f[152]; // c8t368i36
	assign leaf[585] = !f[679] && !f[273] && !f[710] && !f[438]; // c8t378i37
	assign leaf[586] = !f[679] && !f[273] && !f[710] && f[438]; // c8t378i37
	assign leaf[587] = !f[679] && !f[273] && f[710] && !f[542]; // c8t378i37
	assign leaf[588] = !f[679] && !f[273] && f[710] && f[542]; // c8t378i37
	assign leaf[589] = !f[679] && f[273] && !f[480] && !f[243]; // c8t378i37
	assign leaf[590] = !f[679] && f[273] && !f[480] && f[243]; // c8t378i37
	assign leaf[591] = !f[679] && f[273] && f[480] && !f[633]; // c8t378i37
	assign leaf[592] = !f[679] && f[273] && f[480] && f[633]; // c8t378i37
	assign leaf[593] = f[679] && !f[540] && !f[711] && !f[538]; // c8t378i37
	assign leaf[594] = f[679] && !f[540] && !f[711] && f[538]; // c8t378i37
	assign leaf[595] = f[679] && !f[540] && f[711] && !f[182]; // c8t378i37
	assign leaf[596] = f[679] && !f[540] && f[711] && f[182]; // c8t378i37
	assign leaf[597] = f[679] && f[540] && !f[681] && !f[621]; // c8t378i37
	assign leaf[598] = f[679] && f[540] && !f[681] && f[621]; // c8t378i37
	assign leaf[599] = f[679] && f[540] && f[681] && !f[232]; // c8t378i37
	assign leaf[600] = f[679] && f[540] && f[681] && f[232]; // c8t378i37
	assign leaf[601] = !f[399] && !f[317] && !f[292] && !f[265]; // c8t388i38
	assign leaf[602] = !f[399] && !f[317] && !f[292] && f[265]; // c8t388i38
	assign leaf[603] = !f[399] && !f[317] && f[292] && !f[347]; // c8t388i38
	assign leaf[604] = !f[399] && !f[317] && f[292] && f[347]; // c8t388i38
	assign leaf[605] = !f[399] && f[317] && !f[290] && !f[372]; // c8t388i38
	assign leaf[606] = !f[399] && f[317] && !f[290] && f[372]; // c8t388i38
	assign leaf[607] = !f[399] && f[317] && f[290] && !f[517]; // c8t388i38
	assign leaf[608] = !f[399] && f[317] && f[290] && f[517]; // c8t388i38
	assign leaf[609] = f[399] && !f[607] && !f[304] && !f[287]; // c8t388i38
	assign leaf[610] = f[399] && !f[607] && !f[304] && f[287]; // c8t388i38
	assign leaf[611] = f[399] && !f[607] && f[304] && !f[212]; // c8t388i38
	assign leaf[612] = f[399] && !f[607] && f[304] && f[212]; // c8t388i38
	assign leaf[613] = f[399] && f[607] && !f[489] && !f[523]; // c8t388i38
	assign leaf[614] = f[399] && f[607] && !f[489] && f[523]; // c8t388i38
	assign leaf[615] = f[399] && f[607] && f[489] && !f[374]; // c8t388i38
	assign leaf[616] = f[399] && f[607] && f[489] && f[374]; // c8t388i38
	assign leaf[617] = !f[219] && !f[412] && !f[688] && !f[350]; // c8t398i39
	assign leaf[618] = !f[219] && !f[412] && !f[688] && f[350]; // c8t398i39
	assign leaf[619] = !f[219] && !f[412] && f[688] && !f[545]; // c8t398i39
	assign leaf[620] = !f[219] && !f[412] && f[688] && f[545]; // c8t398i39
	assign leaf[621] = !f[219] && f[412] && !f[332] && !f[126]; // c8t398i39
	assign leaf[622] = !f[219] && f[412] && !f[332] && f[126]; // c8t398i39
	assign leaf[623] = !f[219] && f[412] && f[332] && !f[344]; // c8t398i39
	assign leaf[624] = !f[219] && f[412] && f[332] && f[344]; // c8t398i39
	assign leaf[625] = f[219] && !f[454] && !f[649] && !f[379]; // c8t398i39
	assign leaf[626] = f[219] && !f[454] && !f[649] && f[379]; // c8t398i39
	assign leaf[627] = f[219] && !f[454] && f[649] && !f[597]; // c8t398i39
	assign leaf[628] = f[219] && !f[454] && f[649] && f[597]; // c8t398i39
	assign leaf[629] = f[219] && f[454] && !f[272] && !f[181]; // c8t398i39
	assign leaf[630] = f[219] && f[454] && !f[272] && f[181]; // c8t398i39
	assign leaf[631] = f[219] && f[454] && f[272] && !f[595]; // c8t398i39
	assign leaf[632] = f[219] && f[454] && f[272] && f[595]; // c8t398i39
	assign leaf[633] = !f[340] && !f[468] && !f[357] && !f[410]; // c8t408i40
	assign leaf[634] = !f[340] && !f[468] && !f[357] && f[410]; // c8t408i40
	assign leaf[635] = !f[340] && !f[468] && f[357] && !f[326]; // c8t408i40
	assign leaf[636] = !f[340] && !f[468] && f[357] && f[326]; // c8t408i40
	assign leaf[637] = !f[340] && f[468] && !f[577] && !f[492]; // c8t408i40
	assign leaf[638] = !f[340] && f[468] && !f[577] && f[492]; // c8t408i40
	assign leaf[639] = !f[340] && f[468] && f[577] && !f[380]; // c8t408i40
	assign leaf[640] = !f[340] && f[468] && f[577] && f[380]; // c8t408i40
	assign leaf[641] = f[340] && !f[464]; // c8t408i40
	assign leaf[642] = f[340] && f[464] && !f[152] && !f[321]; // c8t408i40
	assign leaf[643] = f[340] && f[464] && !f[152] && f[321]; // c8t408i40
	assign leaf[644] = f[340] && f[464] && f[152]; // c8t408i40
	assign leaf[645] = !f[437] && !f[492] && !f[547] && !f[543]; // c8t418i41
	assign leaf[646] = !f[437] && !f[492] && !f[547] && f[543]; // c8t418i41
	assign leaf[647] = !f[437] && !f[492] && f[547] && !f[550]; // c8t418i41
	assign leaf[648] = !f[437] && !f[492] && f[547] && f[550]; // c8t418i41
	assign leaf[649] = !f[437] && f[492] && !f[406] && !f[219]; // c8t418i41
	assign leaf[650] = !f[437] && f[492] && !f[406] && f[219]; // c8t418i41
	assign leaf[651] = !f[437] && f[492] && f[406] && !f[518]; // c8t418i41
	assign leaf[652] = !f[437] && f[492] && f[406] && f[518]; // c8t418i41
	assign leaf[653] = f[437] && !f[353] && !f[489] && !f[323]; // c8t418i41
	assign leaf[654] = f[437] && !f[353] && !f[489] && f[323]; // c8t418i41
	assign leaf[655] = f[437] && !f[353] && f[489] && !f[483]; // c8t418i41
	assign leaf[656] = f[437] && !f[353] && f[489] && f[483]; // c8t418i41
	assign leaf[657] = f[437] && f[353] && !f[491] && !f[483]; // c8t418i41
	assign leaf[658] = f[437] && f[353] && !f[491] && f[483]; // c8t418i41
	assign leaf[659] = f[437] && f[353] && f[491] && !f[662]; // c8t418i41
	assign leaf[660] = f[437] && f[353] && f[491] && f[662]; // c8t418i41
	assign leaf[661] = !f[303] && !f[650] && !f[244] && !f[637]; // c8t428i42
	assign leaf[662] = !f[303] && !f[650] && !f[244] && f[637]; // c8t428i42
	assign leaf[663] = !f[303] && !f[650] && f[244] && !f[242]; // c8t428i42
	assign leaf[664] = !f[303] && !f[650] && f[244] && f[242]; // c8t428i42
	assign leaf[665] = !f[303] && f[650] && !f[539] && !f[541]; // c8t428i42
	assign leaf[666] = !f[303] && f[650] && !f[539] && f[541]; // c8t428i42
	assign leaf[667] = !f[303] && f[650] && f[539] && !f[634]; // c8t428i42
	assign leaf[668] = !f[303] && f[650] && f[539] && f[634]; // c8t428i42
	assign leaf[669] = f[303] && !f[485] && !f[577] && !f[301]; // c8t428i42
	assign leaf[670] = f[303] && !f[485] && !f[577] && f[301]; // c8t428i42
	assign leaf[671] = f[303] && !f[485] && f[577] && !f[409]; // c8t428i42
	assign leaf[672] = f[303] && !f[485] && f[577] && f[409]; // c8t428i42
	assign leaf[673] = f[303] && f[485] && !f[207] && !f[492]; // c8t428i42
	assign leaf[674] = f[303] && f[485] && !f[207] && f[492]; // c8t428i42
	assign leaf[675] = f[303] && f[485] && f[207] && !f[354]; // c8t428i42
	assign leaf[676] = f[303] && f[485] && f[207] && f[354]; // c8t428i42
	assign leaf[677] = !f[542] && !f[512] && !f[544] && !f[510]; // c8t438i43
	assign leaf[678] = !f[542] && !f[512] && !f[544] && f[510]; // c8t438i43
	assign leaf[679] = !f[542] && !f[512] && f[544] && !f[549]; // c8t438i43
	assign leaf[680] = !f[542] && !f[512] && f[544] && f[549]; // c8t438i43
	assign leaf[681] = !f[542] && f[512] && !f[322] && !f[403]; // c8t438i43
	assign leaf[682] = !f[542] && f[512] && !f[322] && f[403]; // c8t438i43
	assign leaf[683] = !f[542] && f[512] && f[322] && !f[540]; // c8t438i43
	assign leaf[684] = !f[542] && f[512] && f[322] && f[540]; // c8t438i43
	assign leaf[685] = f[542] && !f[511] && !f[544] && !f[518]; // c8t438i43
	assign leaf[686] = f[542] && !f[511] && !f[544] && f[518]; // c8t438i43
	assign leaf[687] = f[542] && !f[511] && f[544] && !f[296]; // c8t438i43
	assign leaf[688] = f[542] && !f[511] && f[544] && f[296]; // c8t438i43
	assign leaf[689] = f[542] && f[511] && !f[681] && !f[634]; // c8t438i43
	assign leaf[690] = f[542] && f[511] && !f[681] && f[634]; // c8t438i43
	assign leaf[691] = f[542] && f[511] && f[681] && !f[491]; // c8t438i43
	assign leaf[692] = f[542] && f[511] && f[681] && f[491]; // c8t438i43
	assign leaf[693] = !f[341] && !f[688] && !f[542] && !f[511]; // c8t448i44
	assign leaf[694] = !f[341] && !f[688] && !f[542] && f[511]; // c8t448i44
	assign leaf[695] = !f[341] && !f[688] && f[542] && !f[511]; // c8t448i44
	assign leaf[696] = !f[341] && !f[688] && f[542] && f[511]; // c8t448i44
	assign leaf[697] = !f[341] && f[688] && !f[632] && !f[550]; // c8t448i44
	assign leaf[698] = !f[341] && f[688] && !f[632] && f[550]; // c8t448i44
	assign leaf[699] = !f[341] && f[688] && f[632] && !f[546]; // c8t448i44
	assign leaf[700] = !f[341] && f[688] && f[632] && f[546]; // c8t448i44
	assign leaf[701] = f[341] && !f[315] && !f[636]; // c8t448i44
	assign leaf[702] = f[341] && !f[315] && f[636]; // c8t448i44
	assign leaf[703] = f[341] && f[315] && !f[491] && !f[487]; // c8t448i44
	assign leaf[704] = f[341] && f[315] && !f[491] && f[487]; // c8t448i44
	assign leaf[705] = f[341] && f[315] && f[491] && !f[350]; // c8t448i44
	assign leaf[706] = f[341] && f[315] && f[491] && f[350]; // c8t448i44
	assign leaf[707] = !f[325] && !f[354] && !f[268] && !f[356]; // c8t458i45
	assign leaf[708] = !f[325] && !f[354] && !f[268] && f[356]; // c8t458i45
	assign leaf[709] = !f[325] && !f[354] && f[268] && !f[632]; // c8t458i45
	assign leaf[710] = !f[325] && !f[354] && f[268] && f[632]; // c8t458i45
	assign leaf[711] = !f[325] && f[354] && !f[411] && !f[593]; // c8t458i45
	assign leaf[712] = !f[325] && f[354] && !f[411] && f[593]; // c8t458i45
	assign leaf[713] = !f[325] && f[354] && f[411] && !f[554]; // c8t458i45
	assign leaf[714] = !f[325] && f[354] && f[411] && f[554]; // c8t458i45
	assign leaf[715] = f[325] && !f[409] && !f[492] && !f[518]; // c8t458i45
	assign leaf[716] = f[325] && !f[409] && !f[492] && f[518]; // c8t458i45
	assign leaf[717] = f[325] && !f[409] && f[492] && !f[403]; // c8t458i45
	assign leaf[718] = f[325] && !f[409] && f[492] && f[403]; // c8t458i45
	assign leaf[719] = f[325] && f[409] && !f[495] && !f[351]; // c8t458i45
	assign leaf[720] = f[325] && f[409] && !f[495] && f[351]; // c8t458i45
	assign leaf[721] = f[325] && f[409] && f[495] && !f[426]; // c8t458i45
	assign leaf[722] = f[325] && f[409] && f[495] && f[426]; // c8t458i45
	assign leaf[723] = !f[649] && !f[201] && !f[663] && !f[494]; // c8t468i46
	assign leaf[724] = !f[649] && !f[201] && !f[663] && f[494]; // c8t468i46
	assign leaf[725] = !f[649] && !f[201] && f[663] && !f[574]; // c8t468i46
	assign leaf[726] = !f[649] && !f[201] && f[663] && f[574]; // c8t468i46
	assign leaf[727] = !f[649] && f[201] && !f[318] && !f[342]; // c8t468i46
	assign leaf[728] = !f[649] && f[201] && !f[318] && f[342]; // c8t468i46
	assign leaf[729] = !f[649] && f[201] && f[318] && !f[296]; // c8t468i46
	assign leaf[730] = !f[649] && f[201] && f[318] && f[296]; // c8t468i46
	assign leaf[731] = f[649] && !f[624] && !f[568]; // c8t468i46
	assign leaf[732] = f[649] && !f[624] && f[568]; // c8t468i46
	assign leaf[733] = f[649] && f[624] && !f[456] && !f[348]; // c8t468i46
	assign leaf[734] = f[649] && f[624] && !f[456] && f[348]; // c8t468i46
	assign leaf[735] = f[649] && f[624] && f[456] && !f[437]; // c8t468i46
	assign leaf[736] = f[649] && f[624] && f[456] && f[437]; // c8t468i46
	assign leaf[737] = !f[238] && !f[321] && !f[347] && !f[374]; // c8t478i47
	assign leaf[738] = !f[238] && !f[321] && !f[347] && f[374]; // c8t478i47
	assign leaf[739] = !f[238] && !f[321] && f[347] && !f[402]; // c8t478i47
	assign leaf[740] = !f[238] && !f[321] && f[347] && f[402]; // c8t478i47
	assign leaf[741] = !f[238] && f[321] && !f[346] && !f[154]; // c8t478i47
	assign leaf[742] = !f[238] && f[321] && !f[346] && f[154]; // c8t478i47
	assign leaf[743] = !f[238] && f[321] && f[346] && !f[456]; // c8t478i47
	assign leaf[744] = !f[238] && f[321] && f[346] && f[456]; // c8t478i47
	assign leaf[745] = f[238] && !f[304] && !f[188] && !f[663]; // c8t478i47
	assign leaf[746] = f[238] && !f[304] && !f[188] && f[663]; // c8t478i47
	assign leaf[747] = f[238] && !f[304] && f[188] && !f[633]; // c8t478i47
	assign leaf[748] = f[238] && !f[304] && f[188] && f[633]; // c8t478i47
	assign leaf[749] = f[238] && f[304] && !f[400] && !f[520]; // c8t478i47
	assign leaf[750] = f[238] && f[304] && !f[400] && f[520]; // c8t478i47
	assign leaf[751] = f[238] && f[304] && f[400] && !f[348]; // c8t478i47
	assign leaf[752] = f[238] && f[304] && f[400] && f[348]; // c8t478i47
	assign leaf[753] = !f[273] && !f[289] && !f[375] && !f[320]; // c8t488i48
	assign leaf[754] = !f[273] && !f[289] && !f[375] && f[320]; // c8t488i48
	assign leaf[755] = !f[273] && !f[289] && f[375] && !f[315]; // c8t488i48
	assign leaf[756] = !f[273] && !f[289] && f[375] && f[315]; // c8t488i48
	assign leaf[757] = !f[273] && f[289] && !f[375] && !f[320]; // c8t488i48
	assign leaf[758] = !f[273] && f[289] && !f[375] && f[320]; // c8t488i48
	assign leaf[759] = !f[273] && f[289] && f[375] && !f[401]; // c8t488i48
	assign leaf[760] = !f[273] && f[289] && f[375] && f[401]; // c8t488i48
	assign leaf[761] = f[273] && !f[322] && !f[402] && !f[348]; // c8t488i48
	assign leaf[762] = f[273] && !f[322] && !f[402] && f[348]; // c8t488i48
	assign leaf[763] = f[273] && !f[322] && f[402] && !f[288]; // c8t488i48
	assign leaf[764] = f[273] && !f[322] && f[402] && f[288]; // c8t488i48
	assign leaf[765] = f[273] && f[322] && !f[347] && !f[261]; // c8t488i48
	assign leaf[766] = f[273] && f[322] && !f[347] && f[261]; // c8t488i48
	assign leaf[767] = f[273] && f[322] && f[347] && !f[519]; // c8t488i48
	assign leaf[768] = f[273] && f[322] && f[347] && f[519]; // c8t488i48
	assign leaf[769] = !f[441] && !f[678] && !f[289] && !f[375]; // c8t498i49
	assign leaf[770] = !f[441] && !f[678] && !f[289] && f[375]; // c8t498i49
	assign leaf[771] = !f[441] && !f[678] && f[289] && !f[545]; // c8t498i49
	assign leaf[772] = !f[441] && !f[678] && f[289] && f[545]; // c8t498i49
	assign leaf[773] = !f[441] && f[678] && !f[512] && !f[406]; // c8t498i49
	assign leaf[774] = !f[441] && f[678] && !f[512] && f[406]; // c8t498i49
	assign leaf[775] = !f[441] && f[678] && f[512] && !f[566]; // c8t498i49
	assign leaf[776] = !f[441] && f[678] && f[512] && f[566]; // c8t498i49
	assign leaf[777] = f[441] && !f[523] && !f[411] && !f[596]; // c8t498i49
	assign leaf[778] = f[441] && !f[523] && !f[411] && f[596]; // c8t498i49
	assign leaf[779] = f[441] && !f[523] && f[411] && !f[160]; // c8t498i49
	assign leaf[780] = f[441] && !f[523] && f[411] && f[160]; // c8t498i49
	assign leaf[781] = f[441] && f[523] && !f[218] && !f[214]; // c8t498i49
	assign leaf[782] = f[441] && f[523] && !f[218] && f[214]; // c8t498i49
	assign leaf[783] = f[441] && f[523] && f[218] && !f[239]; // c8t498i49
	assign leaf[784] = f[441] && f[523] && f[218] && f[239]; // c8t498i49
	assign leaf[785] = !f[705] && !f[219] && !f[708] && !f[120]; // c8t508i50
	assign leaf[786] = !f[705] && !f[219] && !f[708] && f[120]; // c8t508i50
	assign leaf[787] = !f[705] && !f[219] && f[708] && !f[568]; // c8t508i50
	assign leaf[788] = !f[705] && !f[219] && f[708] && f[568]; // c8t508i50
	assign leaf[789] = !f[705] && f[219] && !f[379] && !f[543]; // c8t508i50
	assign leaf[790] = !f[705] && f[219] && !f[379] && f[543]; // c8t508i50
	assign leaf[791] = !f[705] && f[219] && f[379] && !f[346]; // c8t508i50
	assign leaf[792] = !f[705] && f[219] && f[379] && f[346]; // c8t508i50
	assign leaf[793] = f[705]; // c8t508i50
	assign leaf[794] = !f[452] && !f[333] && !f[705] && !f[563]; // c8t518i51
	assign leaf[795] = !f[452] && !f[333] && !f[705] && f[563]; // c8t518i51
	assign leaf[796] = !f[452] && !f[333] && f[705]; // c8t518i51
	assign leaf[797] = !f[452] && f[333] && !f[299] && !f[573]; // c8t518i51
	assign leaf[798] = !f[452] && f[333] && !f[299] && f[573]; // c8t518i51
	assign leaf[799] = !f[452] && f[333] && f[299]; // c8t518i51
	assign leaf[800] = f[452]; // c8t518i51
	assign leaf[801] = !f[304] && !f[708] && !f[322] && !f[462]; // c8t528i52
	assign leaf[802] = !f[304] && !f[708] && !f[322] && f[462]; // c8t528i52
	assign leaf[803] = !f[304] && !f[708] && f[322] && !f[546]; // c8t528i52
	assign leaf[804] = !f[304] && !f[708] && f[322] && f[546]; // c8t528i52
	assign leaf[805] = !f[304] && f[708] && !f[568] && !f[630]; // c8t528i52
	assign leaf[806] = !f[304] && f[708] && !f[568] && f[630]; // c8t528i52
	assign leaf[807] = !f[304] && f[708] && f[568]; // c8t528i52
	assign leaf[808] = f[304] && !f[322] && !f[486] && !f[653]; // c8t528i52
	assign leaf[809] = f[304] && !f[322] && !f[486] && f[653]; // c8t528i52
	assign leaf[810] = f[304] && !f[322] && f[486]; // c8t528i52
	assign leaf[811] = f[304] && f[322] && !f[212] && !f[268]; // c8t528i52
	assign leaf[812] = f[304] && f[322] && !f[212] && f[268]; // c8t528i52
	assign leaf[813] = f[304] && f[322] && f[212] && !f[262]; // c8t528i52
	assign leaf[814] = f[304] && f[322] && f[212] && f[262]; // c8t528i52
	assign leaf[815] = !f[649] && !f[708] && !f[434] && !f[429]; // c8t538i53
	assign leaf[816] = !f[649] && !f[708] && !f[434] && f[429]; // c8t538i53
	assign leaf[817] = !f[649] && !f[708] && f[434] && !f[100]; // c8t538i53
	assign leaf[818] = !f[649] && !f[708] && f[434] && f[100]; // c8t538i53
	assign leaf[819] = !f[649] && f[708] && !f[513] && !f[575]; // c8t538i53
	assign leaf[820] = !f[649] && f[708] && !f[513] && f[575]; // c8t538i53
	assign leaf[821] = !f[649] && f[708] && f[513]; // c8t538i53
	assign leaf[822] = f[649] && !f[539] && !f[247]; // c8t538i53
	assign leaf[823] = f[649] && !f[539] && f[247]; // c8t538i53
	assign leaf[824] = f[649] && f[539] && !f[347] && !f[349]; // c8t538i53
	assign leaf[825] = f[649] && f[539] && !f[347] && f[349]; // c8t538i53
	assign leaf[826] = f[649] && f[539] && f[347]; // c8t538i53
	assign leaf[827] = !f[176] && !f[687] && !f[630] && !f[575]; // c8t548i54
	assign leaf[828] = !f[176] && !f[687] && !f[630] && f[575]; // c8t548i54
	assign leaf[829] = !f[176] && !f[687] && f[630] && !f[657]; // c8t548i54
	assign leaf[830] = !f[176] && !f[687] && f[630] && f[657]; // c8t548i54
	assign leaf[831] = !f[176] && f[687] && !f[631] && !f[689]; // c8t548i54
	assign leaf[832] = !f[176] && f[687] && !f[631] && f[689]; // c8t548i54
	assign leaf[833] = !f[176] && f[687] && f[631] && !f[545]; // c8t548i54
	assign leaf[834] = !f[176] && f[687] && f[631] && f[545]; // c8t548i54
	assign leaf[835] = f[176] && !f[657] && !f[636] && !f[628]; // c8t548i54
	assign leaf[836] = f[176] && !f[657] && !f[636] && f[628]; // c8t548i54
	assign leaf[837] = f[176] && !f[657] && f[636] && !f[631]; // c8t548i54
	assign leaf[838] = f[176] && !f[657] && f[636] && f[631]; // c8t548i54
	assign leaf[839] = f[176] && f[657] && !f[209] && !f[128]; // c8t548i54
	assign leaf[840] = f[176] && f[657] && !f[209] && f[128]; // c8t548i54
	assign leaf[841] = f[176] && f[657] && f[209] && !f[492]; // c8t548i54
	assign leaf[842] = f[176] && f[657] && f[209] && f[492]; // c8t548i54
	assign leaf[843] = !f[525] && !f[570] && !f[540] && !f[572]; // c8t558i55
	assign leaf[844] = !f[525] && !f[570] && !f[540] && f[572]; // c8t558i55
	assign leaf[845] = !f[525] && !f[570] && f[540] && !f[604]; // c8t558i55
	assign leaf[846] = !f[525] && !f[570] && f[540] && f[604]; // c8t558i55
	assign leaf[847] = !f[525] && f[570] && !f[572] && !f[518]; // c8t558i55
	assign leaf[848] = !f[525] && f[570] && !f[572] && f[518]; // c8t558i55
	assign leaf[849] = !f[525] && f[570] && f[572] && !f[296]; // c8t558i55
	assign leaf[850] = !f[525] && f[570] && f[572] && f[296]; // c8t558i55
	assign leaf[851] = f[525] && !f[470] && !f[296] && !f[523]; // c8t558i55
	assign leaf[852] = f[525] && !f[470] && !f[296] && f[523]; // c8t558i55
	assign leaf[853] = f[525] && !f[470] && f[296] && !f[550]; // c8t558i55
	assign leaf[854] = f[525] && !f[470] && f[296] && f[550]; // c8t558i55
	assign leaf[855] = f[525] && f[470] && !f[456] && !f[438]; // c8t558i55
	assign leaf[856] = f[525] && f[470] && !f[456] && f[438]; // c8t558i55
	assign leaf[857] = f[525] && f[470] && f[456] && !f[125]; // c8t558i55
	assign leaf[858] = f[525] && f[470] && f[456] && f[125]; // c8t558i55
	assign leaf[859] = !f[341] && !f[277] && !f[679] && !f[302]; // c8t568i56
	assign leaf[860] = !f[341] && !f[277] && !f[679] && f[302]; // c8t568i56
	assign leaf[861] = !f[341] && !f[277] && f[679] && !f[540]; // c8t568i56
	assign leaf[862] = !f[341] && !f[277] && f[679] && f[540]; // c8t568i56
	assign leaf[863] = !f[341] && f[277] && !f[401]; // c8t568i56
	assign leaf[864] = !f[341] && f[277] && f[401] && !f[383]; // c8t568i56
	assign leaf[865] = !f[341] && f[277] && f[401] && f[383]; // c8t568i56
	assign leaf[866] = f[341] && !f[315] && !f[625] && !f[177]; // c8t568i56
	assign leaf[867] = f[341] && !f[315] && !f[625] && f[177]; // c8t568i56
	assign leaf[868] = f[341] && !f[315] && f[625]; // c8t568i56
	assign leaf[869] = f[341] && f[315] && !f[264] && !f[572]; // c8t568i56
	assign leaf[870] = f[341] && f[315] && !f[264] && f[572]; // c8t568i56
	assign leaf[871] = f[341] && f[315] && f[264] && !f[383]; // c8t568i56
	assign leaf[872] = f[341] && f[315] && f[264] && f[383]; // c8t568i56
	assign leaf[873] = !f[165] && !f[381] && !f[464] && !f[491]; // c8t578i57
	assign leaf[874] = !f[165] && !f[381] && !f[464] && f[491]; // c8t578i57
	assign leaf[875] = !f[165] && !f[381] && f[464] && !f[376]; // c8t578i57
	assign leaf[876] = !f[165] && !f[381] && f[464] && f[376]; // c8t578i57
	assign leaf[877] = !f[165] && f[381] && !f[297] && !f[295]; // c8t578i57
	assign leaf[878] = !f[165] && f[381] && !f[297] && f[295]; // c8t578i57
	assign leaf[879] = !f[165] && f[381] && f[297] && !f[180]; // c8t578i57
	assign leaf[880] = !f[165] && f[381] && f[297] && f[180]; // c8t578i57
	assign leaf[881] = f[165]; // c8t578i57
	assign leaf[882] = !f[439] && !f[525] && !f[542] && !f[660]; // c8t588i58
	assign leaf[883] = !f[439] && !f[525] && !f[542] && f[660]; // c8t588i58
	assign leaf[884] = !f[439] && !f[525] && f[542] && !f[538]; // c8t588i58
	assign leaf[885] = !f[439] && !f[525] && f[542] && f[538]; // c8t588i58
	assign leaf[886] = !f[439] && f[525] && !f[456] && !f[467]; // c8t588i58
	assign leaf[887] = !f[439] && f[525] && !f[456] && f[467]; // c8t588i58
	assign leaf[888] = !f[439] && f[525] && f[456] && !f[246]; // c8t588i58
	assign leaf[889] = !f[439] && f[525] && f[456] && f[246]; // c8t588i58
	assign leaf[890] = f[439] && !f[154] && !f[354] && !f[572]; // c8t588i58
	assign leaf[891] = f[439] && !f[154] && !f[354] && f[572]; // c8t588i58
	assign leaf[892] = f[439] && !f[154] && f[354] && !f[625]; // c8t588i58
	assign leaf[893] = f[439] && !f[154] && f[354] && f[625]; // c8t588i58
	assign leaf[894] = f[439] && f[154] && !f[318] && !f[265]; // c8t588i58
	assign leaf[895] = f[439] && f[154] && !f[318] && f[265]; // c8t588i58
	assign leaf[896] = f[439] && f[154] && f[318] && !f[379]; // c8t588i58
	assign leaf[897] = f[439] && f[154] && f[318] && f[379]; // c8t588i58
	assign leaf[898] = !f[276] && !f[284] && !f[684] && !f[601]; // c8t598i59
	assign leaf[899] = !f[276] && !f[284] && !f[684] && f[601]; // c8t598i59
	assign leaf[900] = !f[276] && !f[284] && f[684] && !f[601]; // c8t598i59
	assign leaf[901] = !f[276] && !f[284] && f[684] && f[601]; // c8t598i59
	assign leaf[902] = !f[276] && f[284] && !f[374] && !f[354]; // c8t598i59
	assign leaf[903] = !f[276] && f[284] && !f[374] && f[354]; // c8t598i59
	assign leaf[904] = !f[276] && f[284] && f[374]; // c8t598i59
	assign leaf[905] = f[276] && !f[403] && !f[543]; // c8t598i59
	assign leaf[906] = f[276] && !f[403] && f[543] && !f[299]; // c8t598i59
	assign leaf[907] = f[276] && !f[403] && f[543] && f[299]; // c8t598i59
	assign leaf[908] = f[276] && f[403] && !f[207] && !f[511]; // c8t598i59
	assign leaf[909] = f[276] && f[403] && !f[207] && f[511]; // c8t598i59
	assign leaf[910] = f[276] && f[403] && f[207] && !f[682]; // c8t598i59
	assign leaf[911] = f[276] && f[403] && f[207] && f[682]; // c8t598i59
	assign leaf[912] = !f[469] && !f[317] && !f[627] && !f[653]; // c8t608i60
	assign leaf[913] = !f[469] && !f[317] && !f[627] && f[653]; // c8t608i60
	assign leaf[914] = !f[469] && !f[317] && f[627] && !f[600]; // c8t608i60
	assign leaf[915] = !f[469] && !f[317] && f[627] && f[600]; // c8t608i60
	assign leaf[916] = !f[469] && f[317] && !f[375] && !f[430]; // c8t608i60
	assign leaf[917] = !f[469] && f[317] && !f[375] && f[430]; // c8t608i60
	assign leaf[918] = !f[469] && f[317] && f[375] && !f[401]; // c8t608i60
	assign leaf[919] = !f[469] && f[317] && f[375] && f[401]; // c8t608i60
	assign leaf[920] = f[469] && !f[523] && !f[180] && !f[569]; // c8t608i60
	assign leaf[921] = f[469] && !f[523] && !f[180] && f[569]; // c8t608i60
	assign leaf[922] = f[469] && !f[523] && f[180] && !f[314]; // c8t608i60
	assign leaf[923] = f[469] && !f[523] && f[180] && f[314]; // c8t608i60
	assign leaf[924] = f[469] && f[523] && !f[218] && !f[638]; // c8t608i60
	assign leaf[925] = f[469] && f[523] && !f[218] && f[638]; // c8t608i60
	assign leaf[926] = f[469] && f[523] && f[218] && !f[574]; // c8t608i60
	assign leaf[927] = f[469] && f[523] && f[218] && f[574]; // c8t608i60
	assign leaf[928] = !f[466] && !f[549] && !f[575] && !f[324]; // c8t618i61
	assign leaf[929] = !f[466] && !f[549] && !f[575] && f[324]; // c8t618i61
	assign leaf[930] = !f[466] && !f[549] && f[575] && !f[659]; // c8t618i61
	assign leaf[931] = !f[466] && !f[549] && f[575] && f[659]; // c8t618i61
	assign leaf[932] = !f[466] && f[549] && !f[576] && !f[523]; // c8t618i61
	assign leaf[933] = !f[466] && f[549] && !f[576] && f[523]; // c8t618i61
	assign leaf[934] = !f[466] && f[549] && f[576] && !f[178]; // c8t618i61
	assign leaf[935] = !f[466] && f[549] && f[576] && f[178]; // c8t618i61
	assign leaf[936] = f[466] && !f[520] && !f[436] && !f[267]; // c8t618i61
	assign leaf[937] = f[466] && !f[520] && !f[436] && f[267]; // c8t618i61
	assign leaf[938] = f[466] && !f[520] && f[436] && !f[351]; // c8t618i61
	assign leaf[939] = f[466] && !f[520] && f[436] && f[351]; // c8t618i61
	assign leaf[940] = f[466] && f[520] && !f[284] && !f[594]; // c8t618i61
	assign leaf[941] = f[466] && f[520] && !f[284] && f[594]; // c8t618i61
	assign leaf[942] = f[466] && f[520] && f[284]; // c8t618i61
	assign leaf[943] = !f[437] && !f[291] && !f[657] && !f[573]; // c8t628i62
	assign leaf[944] = !f[437] && !f[291] && !f[657] && f[573]; // c8t628i62
	assign leaf[945] = !f[437] && !f[291] && f[657] && !f[517]; // c8t628i62
	assign leaf[946] = !f[437] && !f[291] && f[657] && f[517]; // c8t628i62
	assign leaf[947] = !f[437] && f[291] && !f[520] && !f[300]; // c8t628i62
	assign leaf[948] = !f[437] && f[291] && !f[520] && f[300]; // c8t628i62
	assign leaf[949] = !f[437] && f[291] && f[520] && !f[351]; // c8t628i62
	assign leaf[950] = !f[437] && f[291] && f[520] && f[351]; // c8t628i62
	assign leaf[951] = f[437] && !f[381] && !f[494] && !f[406]; // c8t628i62
	assign leaf[952] = f[437] && !f[381] && !f[494] && f[406]; // c8t628i62
	assign leaf[953] = f[437] && !f[381] && f[494] && !f[351]; // c8t628i62
	assign leaf[954] = f[437] && !f[381] && f[494] && f[351]; // c8t628i62
	assign leaf[955] = f[437] && f[381] && !f[273] && !f[179]; // c8t628i62
	assign leaf[956] = f[437] && f[381] && !f[273] && f[179]; // c8t628i62
	assign leaf[957] = f[437] && f[381] && f[273] && !f[686]; // c8t628i62
	assign leaf[958] = f[437] && f[381] && f[273] && f[686]; // c8t628i62
	assign leaf[959] = !f[328] && !f[271] && !f[269] && !f[385]; // c8t638i63
	assign leaf[960] = !f[328] && !f[271] && !f[269] && f[385]; // c8t638i63
	assign leaf[961] = !f[328] && !f[271] && f[269] && !f[326]; // c8t638i63
	assign leaf[962] = !f[328] && !f[271] && f[269] && f[326]; // c8t638i63
	assign leaf[963] = !f[328] && f[271] && !f[241] && !f[188]; // c8t638i63
	assign leaf[964] = !f[328] && f[271] && !f[241] && f[188]; // c8t638i63
	assign leaf[965] = !f[328] && f[271] && f[241] && !f[539]; // c8t638i63
	assign leaf[966] = !f[328] && f[271] && f[241] && f[539]; // c8t638i63
	assign leaf[967] = f[328] && !f[298] && !f[385] && !f[295]; // c8t638i63
	assign leaf[968] = f[328] && !f[298] && !f[385] && f[295]; // c8t638i63
	assign leaf[969] = f[328] && !f[298] && f[385] && !f[292]; // c8t638i63
	assign leaf[970] = f[328] && !f[298] && f[385] && f[292]; // c8t638i63
	assign leaf[971] = f[328] && f[298] && !f[240] && !f[356]; // c8t638i63
	assign leaf[972] = f[328] && f[298] && !f[240] && f[356]; // c8t638i63
	assign leaf[973] = f[328] && f[298] && f[240] && !f[650]; // c8t638i63
	assign leaf[974] = f[328] && f[298] && f[240] && f[650]; // c8t638i63
	assign leaf[975] = !f[679] && !f[136] && !f[708] && !f[452]; // c8t648i64
	assign leaf[976] = !f[679] && !f[136] && !f[708] && f[452]; // c8t648i64
	assign leaf[977] = !f[679] && !f[136] && f[708]; // c8t648i64
	assign leaf[978] = !f[679] && f[136]; // c8t648i64
	assign leaf[979] = f[679] && !f[540] && !f[710] && !f[247]; // c8t648i64
	assign leaf[980] = f[679] && !f[540] && !f[710] && f[247]; // c8t648i64
	assign leaf[981] = f[679] && !f[540] && f[710]; // c8t648i64
	assign leaf[982] = f[679] && f[540] && !f[373] && !f[548]; // c8t648i64
	assign leaf[983] = f[679] && f[540] && !f[373] && f[548]; // c8t648i64
	assign leaf[984] = f[679] && f[540] && f[373]; // c8t648i64
	assign leaf[985] = !f[341] && !f[491] && !f[294] && !f[303]; // c8t658i65
	assign leaf[986] = !f[341] && !f[491] && !f[294] && f[303]; // c8t658i65
	assign leaf[987] = !f[341] && !f[491] && f[294] && !f[380]; // c8t658i65
	assign leaf[988] = !f[341] && !f[491] && f[294] && f[380]; // c8t658i65
	assign leaf[989] = !f[341] && f[491] && !f[436] && !f[494]; // c8t658i65
	assign leaf[990] = !f[341] && f[491] && !f[436] && f[494]; // c8t658i65
	assign leaf[991] = !f[341] && f[491] && f[436] && !f[352]; // c8t658i65
	assign leaf[992] = !f[341] && f[491] && f[436] && f[352]; // c8t658i65
	assign leaf[993] = f[341] && !f[315] && !f[662]; // c8t658i65
	assign leaf[994] = f[341] && !f[315] && f[662]; // c8t658i65
	assign leaf[995] = f[341] && f[315] && !f[464] && !f[486]; // c8t658i65
	assign leaf[996] = f[341] && f[315] && !f[464] && f[486]; // c8t658i65
	assign leaf[997] = f[341] && f[315] && f[464] && !f[601]; // c8t658i65
	assign leaf[998] = f[341] && f[315] && f[464] && f[601]; // c8t658i65
	assign leaf[999] = !f[465] && !f[520] && !f[207] && !f[627]; // c8t668i66
	assign leaf[1000] = !f[465] && !f[520] && !f[207] && f[627]; // c8t668i66
	assign leaf[1001] = !f[465] && !f[520] && f[207] && !f[600]; // c8t668i66
	assign leaf[1002] = !f[465] && !f[520] && f[207] && f[600]; // c8t668i66
	assign leaf[1003] = !f[465] && f[520] && !f[434] && !f[602]; // c8t668i66
	assign leaf[1004] = !f[465] && f[520] && !f[434] && f[602]; // c8t668i66
	assign leaf[1005] = !f[465] && f[520] && f[434] && !f[235]; // c8t668i66
	assign leaf[1006] = !f[465] && f[520] && f[434] && f[235]; // c8t668i66
	assign leaf[1007] = f[465] && !f[151] && !f[216] && !f[266]; // c8t668i66
	assign leaf[1008] = f[465] && !f[151] && !f[216] && f[266]; // c8t668i66
	assign leaf[1009] = f[465] && !f[151] && f[216] && !f[125]; // c8t668i66
	assign leaf[1010] = f[465] && !f[151] && f[216] && f[125]; // c8t668i66
	assign leaf[1011] = f[465] && f[151] && !f[487] && !f[313]; // c8t668i66
	assign leaf[1012] = f[465] && f[151] && !f[487] && f[313]; // c8t668i66
	assign leaf[1013] = f[465] && f[151] && f[487] && !f[543]; // c8t668i66
	assign leaf[1014] = f[465] && f[151] && f[487] && f[543]; // c8t668i66
	assign leaf[1015] = !f[382] && !f[326] && !f[263] && !f[290]; // c8t678i67
	assign leaf[1016] = !f[382] && !f[326] && !f[263] && f[290]; // c8t678i67
	assign leaf[1017] = !f[382] && !f[326] && f[263] && !f[296]; // c8t678i67
	assign leaf[1018] = !f[382] && !f[326] && f[263] && f[296]; // c8t678i67
	assign leaf[1019] = !f[382] && f[326] && !f[215] && !f[356]; // c8t678i67
	assign leaf[1020] = !f[382] && f[326] && !f[215] && f[356]; // c8t678i67
	assign leaf[1021] = !f[382] && f[326] && f[215] && !f[296]; // c8t678i67
	assign leaf[1022] = !f[382] && f[326] && f[215] && f[296]; // c8t678i67
	assign leaf[1023] = f[382] && !f[352] && !f[494] && !f[685]; // c8t678i67
	assign leaf[1024] = f[382] && !f[352] && !f[494] && f[685]; // c8t678i67
	assign leaf[1025] = f[382] && !f[352] && f[494] && !f[411]; // c8t678i67
	assign leaf[1026] = f[382] && !f[352] && f[494] && f[411]; // c8t678i67
	assign leaf[1027] = f[382] && f[352] && !f[483] && !f[513]; // c8t678i67
	assign leaf[1028] = f[382] && f[352] && !f[483] && f[513]; // c8t678i67
	assign leaf[1029] = f[382] && f[352] && f[483] && !f[625]; // c8t678i67
	assign leaf[1030] = f[382] && f[352] && f[483] && f[625]; // c8t678i67
	assign leaf[1031] = !f[314] && !f[290] && !f[316] && !f[232]; // c8t688i68
	assign leaf[1032] = !f[314] && !f[290] && !f[316] && f[232]; // c8t688i68
	assign leaf[1033] = !f[314] && !f[290] && f[316] && !f[234]; // c8t688i68
	assign leaf[1034] = !f[314] && !f[290] && f[316] && f[234]; // c8t688i68
	assign leaf[1035] = !f[314] && f[290] && !f[348] && !f[544]; // c8t688i68
	assign leaf[1036] = !f[314] && f[290] && !f[348] && f[544]; // c8t688i68
	assign leaf[1037] = !f[314] && f[290] && f[348] && !f[373]; // c8t688i68
	assign leaf[1038] = !f[314] && f[290] && f[348] && f[373]; // c8t688i68
	assign leaf[1039] = f[314] && !f[353] && !f[373] && !f[495]; // c8t688i68
	assign leaf[1040] = f[314] && !f[353] && !f[373] && f[495]; // c8t688i68
	assign leaf[1041] = f[314] && !f[353] && f[373] && !f[544]; // c8t688i68
	assign leaf[1042] = f[314] && !f[353] && f[373] && f[544]; // c8t688i68
	assign leaf[1043] = f[314] && f[353] && !f[681] && !f[433]; // c8t688i68
	assign leaf[1044] = f[314] && f[353] && !f[681] && f[433]; // c8t688i68
	assign leaf[1045] = f[314] && f[353] && f[681]; // c8t688i68
	assign leaf[1046] = !f[627] && !f[634] && !f[682] && !f[572]; // c8t698i69
	assign leaf[1047] = !f[627] && !f[634] && !f[682] && f[572]; // c8t698i69
	assign leaf[1048] = !f[627] && !f[634] && f[682] && !f[521]; // c8t698i69
	assign leaf[1049] = !f[627] && !f[634] && f[682] && f[521]; // c8t698i69
	assign leaf[1050] = !f[627] && f[634] && !f[574] && !f[601]; // c8t698i69
	assign leaf[1051] = !f[627] && f[634] && !f[574] && f[601]; // c8t698i69
	assign leaf[1052] = !f[627] && f[634] && f[574] && !f[512]; // c8t698i69
	assign leaf[1053] = !f[627] && f[634] && f[574] && f[512]; // c8t698i69
	assign leaf[1054] = f[627] && !f[654] && !f[635] && !f[687]; // c8t698i69
	assign leaf[1055] = f[627] && !f[654] && !f[635] && f[687]; // c8t698i69
	assign leaf[1056] = f[627] && !f[654] && f[635] && !f[207]; // c8t698i69
	assign leaf[1057] = f[627] && !f[654] && f[635] && f[207]; // c8t698i69
	assign leaf[1058] = f[627] && f[654] && !f[600] && !f[293]; // c8t698i69
	assign leaf[1059] = f[627] && f[654] && !f[600] && f[293]; // c8t698i69
	assign leaf[1060] = f[627] && f[654] && f[600] && !f[623]; // c8t698i69
	assign leaf[1061] = f[627] && f[654] && f[600] && f[623]; // c8t698i69
	assign leaf[1062] = !f[682] && !f[627] && !f[633] && !f[689]; // c8t708i70
	assign leaf[1063] = !f[682] && !f[627] && !f[633] && f[689]; // c8t708i70
	assign leaf[1064] = !f[682] && !f[627] && f[633] && !f[513]; // c8t708i70
	assign leaf[1065] = !f[682] && !f[627] && f[633] && f[513]; // c8t708i70
	assign leaf[1066] = !f[682] && f[627] && !f[632] && !f[572]; // c8t708i70
	assign leaf[1067] = !f[682] && f[627] && !f[632] && f[572]; // c8t708i70
	assign leaf[1068] = !f[682] && f[627] && f[632] && !f[601]; // c8t708i70
	assign leaf[1069] = !f[682] && f[627] && f[632] && f[601]; // c8t708i70
	assign leaf[1070] = f[682] && !f[542] && !f[539] && !f[540]; // c8t708i70
	assign leaf[1071] = f[682] && !f[542] && !f[539] && f[540]; // c8t708i70
	assign leaf[1072] = f[682] && !f[542] && f[539] && !f[494]; // c8t708i70
	assign leaf[1073] = f[682] && !f[542] && f[539] && f[494]; // c8t708i70
	assign leaf[1074] = f[682] && f[542] && !f[661] && !f[405]; // c8t708i70
	assign leaf[1075] = f[682] && f[542] && !f[661] && f[405]; // c8t708i70
	assign leaf[1076] = f[682] && f[542] && f[661] && !f[657]; // c8t708i70
	assign leaf[1077] = f[682] && f[542] && f[661] && f[657]; // c8t708i70
	assign leaf[1078] = !f[542] && !f[512] && !f[653] && !f[545]; // c8t718i71
	assign leaf[1079] = !f[542] && !f[512] && !f[653] && f[545]; // c8t718i71
	assign leaf[1080] = !f[542] && !f[512] && f[653] && !f[509]; // c8t718i71
	assign leaf[1081] = !f[542] && !f[512] && f[653] && f[509]; // c8t718i71
	assign leaf[1082] = !f[542] && f[512] && !f[379] && !f[635]; // c8t718i71
	assign leaf[1083] = !f[542] && f[512] && !f[379] && f[635]; // c8t718i71
	assign leaf[1084] = !f[542] && f[512] && f[379] && !f[604]; // c8t718i71
	assign leaf[1085] = !f[542] && f[512] && f[379] && f[604]; // c8t718i71
	assign leaf[1086] = f[542] && !f[512] && !f[324] && !f[576]; // c8t718i71
	assign leaf[1087] = f[542] && !f[512] && !f[324] && f[576]; // c8t718i71
	assign leaf[1088] = f[542] && !f[512] && f[324] && !f[241]; // c8t718i71
	assign leaf[1089] = f[542] && !f[512] && f[324] && f[241]; // c8t718i71
	assign leaf[1090] = f[542] && f[512] && !f[458] && !f[576]; // c8t718i71
	assign leaf[1091] = f[542] && f[512] && !f[458] && f[576]; // c8t718i71
	assign leaf[1092] = f[542] && f[512] && f[458] && !f[682]; // c8t718i71
	assign leaf[1093] = f[542] && f[512] && f[458] && f[682]; // c8t718i71
	assign leaf[1094] = !f[176] && !f[292] && !f[265] && !f[598]; // c8t728i72
	assign leaf[1095] = !f[176] && !f[292] && !f[265] && f[598]; // c8t728i72
	assign leaf[1096] = !f[176] && !f[292] && f[265] && !f[239]; // c8t728i72
	assign leaf[1097] = !f[176] && !f[292] && f[265] && f[239]; // c8t728i72
	assign leaf[1098] = !f[176] && f[292] && !f[349] && !f[685]; // c8t728i72
	assign leaf[1099] = !f[176] && f[292] && !f[349] && f[685]; // c8t728i72
	assign leaf[1100] = !f[176] && f[292] && f[349] && !f[238]; // c8t728i72
	assign leaf[1101] = !f[176] && f[292] && f[349] && f[238]; // c8t728i72
	assign leaf[1102] = f[176] && !f[657] && !f[631] && !f[183]; // c8t728i72
	assign leaf[1103] = f[176] && !f[657] && !f[631] && f[183]; // c8t728i72
	assign leaf[1104] = f[176] && !f[657] && f[631] && !f[607]; // c8t728i72
	assign leaf[1105] = f[176] && !f[657] && f[631] && f[607]; // c8t728i72
	assign leaf[1106] = f[176] && f[657] && !f[321] && !f[630]; // c8t728i72
	assign leaf[1107] = f[176] && f[657] && !f[321] && f[630]; // c8t728i72
	assign leaf[1108] = f[176] && f[657] && f[321] && !f[346]; // c8t728i72
	assign leaf[1109] = f[176] && f[657] && f[321] && f[346]; // c8t728i72
	assign leaf[1110] = !f[214] && !f[265] && !f[461] && !f[345]; // c8t738i73
	assign leaf[1111] = !f[214] && !f[265] && !f[461] && f[345]; // c8t738i73
	assign leaf[1112] = !f[214] && !f[265] && f[461] && !f[320]; // c8t738i73
	assign leaf[1113] = !f[214] && !f[265] && f[461] && f[320]; // c8t738i73
	assign leaf[1114] = !f[214] && f[265] && !f[320] && !f[570]; // c8t738i73
	assign leaf[1115] = !f[214] && f[265] && !f[320] && f[570]; // c8t738i73
	assign leaf[1116] = !f[214] && f[265] && f[320] && !f[162]; // c8t738i73
	assign leaf[1117] = !f[214] && f[265] && f[320] && f[162]; // c8t738i73
	assign leaf[1118] = f[214] && !f[408] && !f[216] && !f[547]; // c8t738i73
	assign leaf[1119] = f[214] && !f[408] && !f[216] && f[547]; // c8t738i73
	assign leaf[1120] = f[214] && !f[408] && f[216] && !f[576]; // c8t738i73
	assign leaf[1121] = f[214] && !f[408] && f[216] && f[576]; // c8t738i73
	assign leaf[1122] = f[214] && f[408] && !f[603] && !f[491]; // c8t738i73
	assign leaf[1123] = f[214] && f[408] && !f[603] && f[491]; // c8t738i73
	assign leaf[1124] = f[214] && f[408] && f[603] && !f[398]; // c8t738i73
	assign leaf[1125] = f[214] && f[408] && f[603] && f[398]; // c8t738i73
	assign leaf[1126] = !f[349] && !f[519] && !f[355] && !f[521]; // c8t748i74
	assign leaf[1127] = !f[349] && !f[519] && !f[355] && f[521]; // c8t748i74
	assign leaf[1128] = !f[349] && !f[519] && f[355] && !f[326]; // c8t748i74
	assign leaf[1129] = !f[349] && !f[519] && f[355] && f[326]; // c8t748i74
	assign leaf[1130] = !f[349] && f[519] && !f[543] && !f[663]; // c8t748i74
	assign leaf[1131] = !f[349] && f[519] && !f[543] && f[663]; // c8t748i74
	assign leaf[1132] = !f[349] && f[519] && f[543] && !f[512]; // c8t748i74
	assign leaf[1133] = !f[349] && f[519] && f[543] && f[512]; // c8t748i74
	assign leaf[1134] = f[349] && !f[519] && !f[436] && !f[544]; // c8t748i74
	assign leaf[1135] = f[349] && !f[519] && !f[436] && f[544]; // c8t748i74
	assign leaf[1136] = f[349] && !f[519] && f[436] && !f[546]; // c8t748i74
	assign leaf[1137] = f[349] && !f[519] && f[436] && f[546]; // c8t748i74
	assign leaf[1138] = f[349] && f[519] && !f[375] && !f[295]; // c8t748i74
	assign leaf[1139] = f[349] && f[519] && !f[375] && f[295]; // c8t748i74
	assign leaf[1140] = f[349] && f[519] && f[375] && !f[579]; // c8t748i74
	assign leaf[1141] = f[349] && f[519] && f[375] && f[579]; // c8t748i74
	assign leaf[1142] = !f[186] && !f[129] && !f[151] && !f[266]; // c8t758i75
	assign leaf[1143] = !f[186] && !f[129] && !f[151] && f[266]; // c8t758i75
	assign leaf[1144] = !f[186] && !f[129] && f[151] && !f[576]; // c8t758i75
	assign leaf[1145] = !f[186] && !f[129] && f[151] && f[576]; // c8t758i75
	assign leaf[1146] = !f[186] && f[129] && !f[378] && !f[517]; // c8t758i75
	assign leaf[1147] = !f[186] && f[129] && !f[378] && f[517]; // c8t758i75
	assign leaf[1148] = !f[186] && f[129] && f[378] && !f[267]; // c8t758i75
	assign leaf[1149] = !f[186] && f[129] && f[378] && f[267]; // c8t758i75
	assign leaf[1150] = f[186] && !f[294] && !f[153] && !f[637]; // c8t758i75
	assign leaf[1151] = f[186] && !f[294] && !f[153] && f[637]; // c8t758i75
	assign leaf[1152] = f[186] && !f[294] && f[153] && !f[599]; // c8t758i75
	assign leaf[1153] = f[186] && !f[294] && f[153] && f[599]; // c8t758i75
	assign leaf[1154] = f[186] && f[294] && !f[348] && !f[319]; // c8t758i75
	assign leaf[1155] = f[186] && f[294] && !f[348] && f[319]; // c8t758i75
	assign leaf[1156] = f[186] && f[294] && f[348] && !f[262]; // c8t758i75
	assign leaf[1157] = f[186] && f[294] && f[348] && f[262]; // c8t758i75
	assign leaf[1158] = !f[236] && !f[260] && !f[262] && !f[238]; // c8t768i76
	assign leaf[1159] = !f[236] && !f[260] && !f[262] && f[238]; // c8t768i76
	assign leaf[1160] = !f[236] && !f[260] && f[262] && !f[240]; // c8t768i76
	assign leaf[1161] = !f[236] && !f[260] && f[262] && f[240]; // c8t768i76
	assign leaf[1162] = !f[236] && f[260] && !f[316] && !f[596]; // c8t768i76
	assign leaf[1163] = !f[236] && f[260] && !f[316] && f[596]; // c8t768i76
	assign leaf[1164] = !f[236] && f[260] && f[316] && !f[271]; // c8t768i76
	assign leaf[1165] = !f[236] && f[260] && f[316] && f[271]; // c8t768i76
	assign leaf[1166] = f[236] && !f[204] && !f[319] && !f[293]; // c8t768i76
	assign leaf[1167] = f[236] && !f[204] && !f[319] && f[293]; // c8t768i76
	assign leaf[1168] = f[236] && !f[204] && f[319] && !f[293]; // c8t768i76
	assign leaf[1169] = f[236] && !f[204] && f[319] && f[293]; // c8t768i76
	assign leaf[1170] = f[236] && f[204] && !f[352] && !f[488]; // c8t768i76
	assign leaf[1171] = f[236] && f[204] && !f[352] && f[488]; // c8t768i76
	assign leaf[1172] = f[236] && f[204] && f[352] && !f[300]; // c8t768i76
	assign leaf[1173] = f[236] && f[204] && f[352] && f[300]; // c8t768i76
	assign leaf[1174] = !f[135] && !f[328] && !f[405] && !f[430]; // c8t778i77
	assign leaf[1175] = !f[135] && !f[328] && !f[405] && f[430]; // c8t778i77
	assign leaf[1176] = !f[135] && !f[328] && f[405] && !f[656]; // c8t778i77
	assign leaf[1177] = !f[135] && !f[328] && f[405] && f[656]; // c8t778i77
	assign leaf[1178] = !f[135] && f[328] && !f[458] && !f[298]; // c8t778i77
	assign leaf[1179] = !f[135] && f[328] && !f[458] && f[298]; // c8t778i77
	assign leaf[1180] = !f[135] && f[328] && f[458] && !f[405]; // c8t778i77
	assign leaf[1181] = !f[135] && f[328] && f[458] && f[405]; // c8t778i77
	assign leaf[1182] = f[135] && !f[270]; // c8t778i77
	assign leaf[1183] = f[135] && f[270]; // c8t778i77
	assign leaf[1184] = !f[508] && !f[399] && !f[276] && !f[549]; // c8t788i78
	assign leaf[1185] = !f[508] && !f[399] && !f[276] && f[549]; // c8t788i78
	assign leaf[1186] = !f[508] && !f[399] && f[276] && !f[298]; // c8t788i78
	assign leaf[1187] = !f[508] && !f[399] && f[276] && f[298]; // c8t788i78
	assign leaf[1188] = !f[508] && f[399] && !f[346] && !f[353]; // c8t788i78
	assign leaf[1189] = !f[508] && f[399] && !f[346] && f[353]; // c8t788i78
	assign leaf[1190] = !f[508] && f[399] && f[346] && !f[432]; // c8t788i78
	assign leaf[1191] = !f[508] && f[399] && f[346] && f[432]; // c8t788i78
	assign leaf[1192] = f[508] && !f[538]; // c8t788i78
	assign leaf[1193] = f[508] && f[538]; // c8t788i78
	assign leaf[1194] = !f[317] && !f[518] && !f[295] && !f[321]; // c8t798i79
	assign leaf[1195] = !f[317] && !f[518] && !f[295] && f[321]; // c8t798i79
	assign leaf[1196] = !f[317] && !f[518] && f[295] && !f[236]; // c8t798i79
	assign leaf[1197] = !f[317] && !f[518] && f[295] && f[236]; // c8t798i79
	assign leaf[1198] = !f[317] && f[518] && !f[597] && !f[372]; // c8t798i79
	assign leaf[1199] = !f[317] && f[518] && !f[597] && f[372]; // c8t798i79
	assign leaf[1200] = !f[317] && f[518] && f[597] && !f[463]; // c8t798i79
	assign leaf[1201] = !f[317] && f[518] && f[597] && f[463]; // c8t798i79
	assign leaf[1202] = f[317] && !f[572] && !f[546] && !f[598]; // c8t798i79
	assign leaf[1203] = f[317] && !f[572] && !f[546] && f[598]; // c8t798i79
	assign leaf[1204] = f[317] && !f[572] && f[546] && !f[606]; // c8t798i79
	assign leaf[1205] = f[317] && !f[572] && f[546] && f[606]; // c8t798i79
	assign leaf[1206] = f[317] && f[572] && !f[685] && !f[431]; // c8t798i79
	assign leaf[1207] = f[317] && f[572] && !f[685] && f[431]; // c8t798i79
	assign leaf[1208] = f[317] && f[572] && f[685] && !f[580]; // c8t798i79
	assign leaf[1209] = f[317] && f[572] && f[685] && f[580]; // c8t798i79
	assign leaf[1210] = !f[408] && !f[181] && !f[371] && !f[353]; // c8t808i80
	assign leaf[1211] = !f[408] && !f[181] && !f[371] && f[353]; // c8t808i80
	assign leaf[1212] = !f[408] && !f[181] && f[371] && !f[216]; // c8t808i80
	assign leaf[1213] = !f[408] && !f[181] && f[371] && f[216]; // c8t808i80
	assign leaf[1214] = !f[408] && f[181] && !f[268] && !f[158]; // c8t808i80
	assign leaf[1215] = !f[408] && f[181] && !f[268] && f[158]; // c8t808i80
	assign leaf[1216] = !f[408] && f[181] && f[268] && !f[602]; // c8t808i80
	assign leaf[1217] = !f[408] && f[181] && f[268] && f[602]; // c8t808i80
	assign leaf[1218] = f[408] && !f[577] && !f[324] && !f[465]; // c8t808i80
	assign leaf[1219] = f[408] && !f[577] && !f[324] && f[465]; // c8t808i80
	assign leaf[1220] = f[408] && !f[577] && f[324] && !f[435]; // c8t808i80
	assign leaf[1221] = f[408] && !f[577] && f[324] && f[435]; // c8t808i80
	assign leaf[1222] = f[408] && f[577] && !f[576] && !f[573]; // c8t808i80
	assign leaf[1223] = f[408] && f[577] && !f[576] && f[573]; // c8t808i80
	assign leaf[1224] = f[408] && f[577] && f[576] && !f[660]; // c8t808i80
	assign leaf[1225] = f[408] && f[577] && f[576] && f[660]; // c8t808i80
	assign leaf[1226] = !f[508] && !f[246] && !f[408] && !f[435]; // c8t818i81
	assign leaf[1227] = !f[508] && !f[246] && !f[408] && f[435]; // c8t818i81
	assign leaf[1228] = !f[508] && !f[246] && f[408] && !f[181]; // c8t818i81
	assign leaf[1229] = !f[508] && !f[246] && f[408] && f[181]; // c8t818i81
	assign leaf[1230] = !f[508] && f[246] && !f[329] && !f[215]; // c8t818i81
	assign leaf[1231] = !f[508] && f[246] && !f[329] && f[215]; // c8t818i81
	assign leaf[1232] = !f[508] && f[246] && f[329] && !f[374]; // c8t818i81
	assign leaf[1233] = !f[508] && f[246] && f[329] && f[374]; // c8t818i81
	assign leaf[1234] = f[508] && !f[153]; // c8t818i81
	assign leaf[1235] = f[508] && f[153]; // c8t818i81
	assign leaf[1236] = !f[302] && !f[235] && !f[234] && !f[348]; // c8t828i82
	assign leaf[1237] = !f[302] && !f[235] && !f[234] && f[348]; // c8t828i82
	assign leaf[1238] = !f[302] && !f[235] && f[234] && !f[291]; // c8t828i82
	assign leaf[1239] = !f[302] && !f[235] && f[234] && f[291]; // c8t828i82
	assign leaf[1240] = !f[302] && f[235] && !f[320] && !f[375]; // c8t828i82
	assign leaf[1241] = !f[302] && f[235] && !f[320] && f[375]; // c8t828i82
	assign leaf[1242] = !f[302] && f[235] && f[320] && !f[349]; // c8t828i82
	assign leaf[1243] = !f[302] && f[235] && f[320] && f[349]; // c8t828i82
	assign leaf[1244] = f[302] && !f[457] && !f[402] && !f[377]; // c8t828i82
	assign leaf[1245] = f[302] && !f[457] && !f[402] && f[377]; // c8t828i82
	assign leaf[1246] = f[302] && !f[457] && f[402] && !f[404]; // c8t828i82
	assign leaf[1247] = f[302] && !f[457] && f[402] && f[404]; // c8t828i82
	assign leaf[1248] = f[302] && f[457] && !f[443] && !f[329]; // c8t828i82
	assign leaf[1249] = f[302] && f[457] && !f[443] && f[329]; // c8t828i82
	assign leaf[1250] = f[302] && f[457] && f[443]; // c8t828i82
	assign leaf[1251] = !f[469] && !f[386] && !f[453] && !f[133]; // c8t838i83
	assign leaf[1252] = !f[469] && !f[386] && !f[453] && f[133]; // c8t838i83
	assign leaf[1253] = !f[469] && !f[386] && f[453]; // c8t838i83
	assign leaf[1254] = !f[469] && f[386] && !f[375] && !f[577]; // c8t838i83
	assign leaf[1255] = !f[469] && f[386] && !f[375] && f[577]; // c8t838i83
	assign leaf[1256] = !f[469] && f[386] && f[375] && !f[300]; // c8t838i83
	assign leaf[1257] = !f[469] && f[386] && f[375] && f[300]; // c8t838i83
	assign leaf[1258] = f[469] && !f[523] && !f[299] && !f[459]; // c8t838i83
	assign leaf[1259] = f[469] && !f[523] && !f[299] && f[459]; // c8t838i83
	assign leaf[1260] = f[469] && !f[523] && f[299] && !f[411]; // c8t838i83
	assign leaf[1261] = f[469] && !f[523] && f[299] && f[411]; // c8t838i83
	assign leaf[1262] = f[469] && f[523] && !f[183] && !f[151]; // c8t838i83
	assign leaf[1263] = f[469] && f[523] && !f[183] && f[151]; // c8t838i83
	assign leaf[1264] = f[469] && f[523] && f[183] && !f[593]; // c8t838i83
	assign leaf[1265] = f[469] && f[523] && f[183] && f[593]; // c8t838i83
	assign leaf[1266] = !f[525] && !f[629] && !f[684] && !f[608]; // c8t848i84
	assign leaf[1267] = !f[525] && !f[629] && !f[684] && f[608]; // c8t848i84
	assign leaf[1268] = !f[525] && !f[629] && f[684] && !f[464]; // c8t848i84
	assign leaf[1269] = !f[525] && !f[629] && f[684] && f[464]; // c8t848i84
	assign leaf[1270] = !f[525] && f[629] && !f[657] && !f[572]; // c8t848i84
	assign leaf[1271] = !f[525] && f[629] && !f[657] && f[572]; // c8t848i84
	assign leaf[1272] = !f[525] && f[629] && f[657] && !f[543]; // c8t848i84
	assign leaf[1273] = !f[525] && f[629] && f[657] && f[543]; // c8t848i84
	assign leaf[1274] = f[525] && !f[458] && !f[571] && !f[522]; // c8t848i84
	assign leaf[1275] = f[525] && !f[458] && !f[571] && f[522]; // c8t848i84
	assign leaf[1276] = f[525] && !f[458] && f[571] && !f[689]; // c8t848i84
	assign leaf[1277] = f[525] && !f[458] && f[571] && f[689]; // c8t848i84
	assign leaf[1278] = f[525] && f[458] && !f[322] && !f[624]; // c8t848i84
	assign leaf[1279] = f[525] && f[458] && !f[322] && f[624]; // c8t848i84
	assign leaf[1280] = f[525] && f[458] && f[322] && !f[385]; // c8t848i84
	assign leaf[1281] = f[525] && f[458] && f[322] && f[385]; // c8t848i84
	assign leaf[1282] = !f[214] && !f[434] && !f[379] && !f[435]; // c8t858i85
	assign leaf[1283] = !f[214] && !f[434] && !f[379] && f[435]; // c8t858i85
	assign leaf[1284] = !f[214] && !f[434] && f[379] && !f[271]; // c8t858i85
	assign leaf[1285] = !f[214] && !f[434] && f[379] && f[271]; // c8t858i85
	assign leaf[1286] = !f[214] && f[434] && !f[293] && !f[348]; // c8t858i85
	assign leaf[1287] = !f[214] && f[434] && !f[293] && f[348]; // c8t858i85
	assign leaf[1288] = !f[214] && f[434] && f[293] && !f[187]; // c8t858i85
	assign leaf[1289] = !f[214] && f[434] && f[293] && f[187]; // c8t858i85
	assign leaf[1290] = f[214] && !f[212] && !f[211] && !f[188]; // c8t858i85
	assign leaf[1291] = f[214] && !f[212] && !f[211] && f[188]; // c8t858i85
	assign leaf[1292] = f[214] && !f[212] && f[211] && !f[239]; // c8t858i85
	assign leaf[1293] = f[214] && !f[212] && f[211] && f[239]; // c8t858i85
	assign leaf[1294] = f[214] && f[212] && !f[329] && !f[482]; // c8t858i85
	assign leaf[1295] = f[214] && f[212] && !f[329] && f[482]; // c8t858i85
	assign leaf[1296] = f[214] && f[212] && f[329] && !f[273]; // c8t858i85
	assign leaf[1297] = f[214] && f[212] && f[329] && f[273]; // c8t858i85
	assign leaf[1298] = !f[125] && !f[439] && !f[525] && !f[592]; // c8t868i86
	assign leaf[1299] = !f[125] && !f[439] && !f[525] && f[592]; // c8t868i86
	assign leaf[1300] = !f[125] && !f[439] && f[525] && !f[187]; // c8t868i86
	assign leaf[1301] = !f[125] && !f[439] && f[525] && f[187]; // c8t868i86
	assign leaf[1302] = !f[125] && f[439] && !f[521] && !f[324]; // c8t868i86
	assign leaf[1303] = !f[125] && f[439] && !f[521] && f[324]; // c8t868i86
	assign leaf[1304] = !f[125] && f[439] && f[521] && !f[303]; // c8t868i86
	assign leaf[1305] = !f[125] && f[439] && f[521] && f[303]; // c8t868i86
	assign leaf[1306] = f[125] && !f[128] && !f[273] && !f[378]; // c8t868i86
	assign leaf[1307] = f[125] && !f[128] && !f[273] && f[378]; // c8t868i86
	assign leaf[1308] = f[125] && !f[128] && f[273]; // c8t868i86
	assign leaf[1309] = f[125] && f[128] && !f[431] && !f[605]; // c8t868i86
	assign leaf[1310] = f[125] && f[128] && !f[431] && f[605]; // c8t868i86
	assign leaf[1311] = f[125] && f[128] && f[431] && !f[296]; // c8t868i86
	assign leaf[1312] = f[125] && f[128] && f[431] && f[296]; // c8t868i86
	assign leaf[1313] = !f[692] && !f[689] && !f[688] && !f[715]; // c8t878i87
	assign leaf[1314] = !f[692] && !f[689] && !f[688] && f[715]; // c8t878i87
	assign leaf[1315] = !f[692] && !f[689] && f[688] && !f[631]; // c8t878i87
	assign leaf[1316] = !f[692] && !f[689] && f[688] && f[631]; // c8t878i87
	assign leaf[1317] = !f[692] && f[689] && !f[493] && !f[631]; // c8t878i87
	assign leaf[1318] = !f[692] && f[689] && !f[493] && f[631]; // c8t878i87
	assign leaf[1319] = !f[692] && f[689] && f[493] && !f[272]; // c8t878i87
	assign leaf[1320] = !f[692] && f[689] && f[493] && f[272]; // c8t878i87
	assign leaf[1321] = f[692] && !f[268] && !f[238]; // c8t878i87
	assign leaf[1322] = f[692] && !f[268] && f[238]; // c8t878i87
	assign leaf[1323] = f[692] && f[268] && !f[575] && !f[460]; // c8t878i87
	assign leaf[1324] = f[692] && f[268] && !f[575] && f[460]; // c8t878i87
	assign leaf[1325] = f[692] && f[268] && f[575]; // c8t878i87
	assign leaf[1326] = !f[678] && !f[161] && !f[570] && !f[632]; // c8t888i88
	assign leaf[1327] = !f[678] && !f[161] && !f[570] && f[632]; // c8t888i88
	assign leaf[1328] = !f[678] && !f[161] && f[570] && !f[572]; // c8t888i88
	assign leaf[1329] = !f[678] && !f[161] && f[570] && f[572]; // c8t888i88
	assign leaf[1330] = !f[678] && f[161] && !f[566] && !f[687]; // c8t888i88
	assign leaf[1331] = !f[678] && f[161] && !f[566] && f[687]; // c8t888i88
	assign leaf[1332] = !f[678] && f[161] && f[566] && !f[569]; // c8t888i88
	assign leaf[1333] = !f[678] && f[161] && f[566] && f[569]; // c8t888i88
	assign leaf[1334] = f[678] && !f[539] && !f[275]; // c8t888i88
	assign leaf[1335] = f[678] && !f[539] && f[275]; // c8t888i88
	assign leaf[1336] = f[678] && f[539]; // c8t888i88
	assign leaf[1337] = !f[149] && !f[603] && !f[605] && !f[540]; // c8t898i89
	assign leaf[1338] = !f[149] && !f[603] && !f[605] && f[540]; // c8t898i89
	assign leaf[1339] = !f[149] && !f[603] && f[605] && !f[689]; // c8t898i89
	assign leaf[1340] = !f[149] && !f[603] && f[605] && f[689]; // c8t898i89
	assign leaf[1341] = !f[149] && f[603] && !f[604] && !f[630]; // c8t898i89
	assign leaf[1342] = !f[149] && f[603] && !f[604] && f[630]; // c8t898i89
	assign leaf[1343] = !f[149] && f[603] && f[604] && !f[427]; // c8t898i89
	assign leaf[1344] = !f[149] && f[603] && f[604] && f[427]; // c8t898i89
	assign leaf[1345] = f[149] && !f[204] && !f[465]; // c8t898i89
	assign leaf[1346] = f[149] && !f[204] && f[465] && !f[293]; // c8t898i89
	assign leaf[1347] = f[149] && !f[204] && f[465] && f[293]; // c8t898i89
	assign leaf[1348] = f[149] && f[204] && !f[319] && !f[239]; // c8t898i89
	assign leaf[1349] = f[149] && f[204] && !f[319] && f[239]; // c8t898i89
	assign leaf[1350] = f[149] && f[204] && f[319] && !f[344]; // c8t898i89
	assign leaf[1351] = f[149] && f[204] && f[319] && f[344]; // c8t898i89
	assign leaf[1352] = !f[486] && !f[488] && !f[517] && !f[456]; // c8t908i90
	assign leaf[1353] = !f[486] && !f[488] && !f[517] && f[456]; // c8t908i90
	assign leaf[1354] = !f[486] && !f[488] && f[517] && !f[549]; // c8t908i90
	assign leaf[1355] = !f[486] && !f[488] && f[517] && f[549]; // c8t908i90
	assign leaf[1356] = !f[486] && f[488] && !f[352] && !f[489]; // c8t908i90
	assign leaf[1357] = !f[486] && f[488] && !f[352] && f[489]; // c8t908i90
	assign leaf[1358] = !f[486] && f[488] && f[352] && !f[290]; // c8t908i90
	assign leaf[1359] = !f[486] && f[488] && f[352] && f[290]; // c8t908i90
	assign leaf[1360] = f[486] && !f[516] && !f[541] && !f[543]; // c8t908i90
	assign leaf[1361] = f[486] && !f[516] && !f[541] && f[543]; // c8t908i90
	assign leaf[1362] = f[486] && !f[516] && f[541] && !f[462]; // c8t908i90
	assign leaf[1363] = f[486] && !f[516] && f[541] && f[462]; // c8t908i90
	assign leaf[1364] = f[486] && f[516] && !f[400] && !f[512]; // c8t908i90
	assign leaf[1365] = f[486] && f[516] && !f[400] && f[512]; // c8t908i90
	assign leaf[1366] = f[486] && f[516] && f[400] && !f[513]; // c8t908i90
	assign leaf[1367] = f[486] && f[516] && f[400] && f[513]; // c8t908i90
	assign leaf[1368] = !f[440] && !f[388] && !f[315] && !f[410]; // c8t918i91
	assign leaf[1369] = !f[440] && !f[388] && !f[315] && f[410]; // c8t918i91
	assign leaf[1370] = !f[440] && !f[388] && f[315] && !f[292]; // c8t918i91
	assign leaf[1371] = !f[440] && !f[388] && f[315] && f[292]; // c8t918i91
	assign leaf[1372] = !f[440] && f[388]; // c8t918i91
	assign leaf[1373] = f[440] && !f[555] && !f[625] && !f[381]; // c8t918i91
	assign leaf[1374] = f[440] && !f[555] && !f[625] && f[381]; // c8t918i91
	assign leaf[1375] = f[440] && !f[555] && f[625] && !f[458]; // c8t918i91
	assign leaf[1376] = f[440] && !f[555] && f[625] && f[458]; // c8t918i91
	assign leaf[1377] = f[440] && f[555] && !f[525]; // c8t918i91
	assign leaf[1378] = f[440] && f[555] && f[525] && !f[354]; // c8t918i91
	assign leaf[1379] = f[440] && f[555] && f[525] && f[354]; // c8t918i91
	assign leaf[1380] = !f[275] && !f[679] && !f[457] && !f[597]; // c8t928i92
	assign leaf[1381] = !f[275] && !f[679] && !f[457] && f[597]; // c8t928i92
	assign leaf[1382] = !f[275] && !f[679] && f[457] && !f[488]; // c8t928i92
	assign leaf[1383] = !f[275] && !f[679] && f[457] && f[488]; // c8t928i92
	assign leaf[1384] = !f[275] && f[679] && !f[540] && !f[378]; // c8t928i92
	assign leaf[1385] = !f[275] && f[679] && !f[540] && f[378]; // c8t928i92
	assign leaf[1386] = !f[275] && f[679] && f[540] && !f[625]; // c8t928i92
	assign leaf[1387] = !f[275] && f[679] && f[540] && f[625]; // c8t928i92
	assign leaf[1388] = f[275] && !f[520] && !f[457] && !f[214]; // c8t928i92
	assign leaf[1389] = f[275] && !f[520] && !f[457] && f[214]; // c8t928i92
	assign leaf[1390] = f[275] && !f[520] && f[457] && !f[485]; // c8t928i92
	assign leaf[1391] = f[275] && !f[520] && f[457] && f[485]; // c8t928i92
	assign leaf[1392] = f[275] && f[520] && !f[207] && !f[466]; // c8t928i92
	assign leaf[1393] = f[275] && f[520] && !f[207] && f[466]; // c8t928i92
	assign leaf[1394] = f[275] && f[520] && f[207] && !f[514]; // c8t928i92
	assign leaf[1395] = f[275] && f[520] && f[207] && f[514]; // c8t928i92
	assign leaf[1396] = !f[341] && !f[214] && !f[601] && !f[656]; // c8t938i93
	assign leaf[1397] = !f[341] && !f[214] && !f[601] && f[656]; // c8t938i93
	assign leaf[1398] = !f[341] && !f[214] && f[601] && !f[656]; // c8t938i93
	assign leaf[1399] = !f[341] && !f[214] && f[601] && f[656]; // c8t938i93
	assign leaf[1400] = !f[341] && f[214] && !f[573] && !f[546]; // c8t938i93
	assign leaf[1401] = !f[341] && f[214] && !f[573] && f[546]; // c8t938i93
	assign leaf[1402] = !f[341] && f[214] && f[573] && !f[435]; // c8t938i93
	assign leaf[1403] = !f[341] && f[214] && f[573] && f[435]; // c8t938i93
	assign leaf[1404] = f[341] && !f[522] && !f[466] && !f[211]; // c8t938i93
	assign leaf[1405] = f[341] && !f[522] && !f[466] && f[211]; // c8t938i93
	assign leaf[1406] = f[341] && !f[522] && f[466]; // c8t938i93
	assign leaf[1407] = f[341] && f[522] && !f[628]; // c8t938i93
	assign leaf[1408] = f[341] && f[522] && f[628]; // c8t938i93
	assign leaf[1409] = !f[657] && !f[629] && !f[381] && !f[317]; // c8t948i94
	assign leaf[1410] = !f[657] && !f[629] && !f[381] && f[317]; // c8t948i94
	assign leaf[1411] = !f[657] && !f[629] && f[381] && !f[433]; // c8t948i94
	assign leaf[1412] = !f[657] && !f[629] && f[381] && f[433]; // c8t948i94
	assign leaf[1413] = !f[657] && f[629] && !f[656] && !f[461]; // c8t948i94
	assign leaf[1414] = !f[657] && f[629] && !f[656] && f[461]; // c8t948i94
	assign leaf[1415] = !f[657] && f[629] && f[656] && !f[492]; // c8t948i94
	assign leaf[1416] = !f[657] && f[629] && f[656] && f[492]; // c8t948i94
	assign leaf[1417] = f[657] && !f[630] && !f[433] && !f[346]; // c8t948i94
	assign leaf[1418] = f[657] && !f[630] && !f[433] && f[346]; // c8t948i94
	assign leaf[1419] = f[657] && !f[630] && f[433] && !f[155]; // c8t948i94
	assign leaf[1420] = f[657] && !f[630] && f[433] && f[155]; // c8t948i94
	assign leaf[1421] = f[657] && f[630] && !f[633] && !f[543]; // c8t948i94
	assign leaf[1422] = f[657] && f[630] && !f[633] && f[543]; // c8t948i94
	assign leaf[1423] = f[657] && f[630] && f[633] && !f[349]; // c8t948i94
	assign leaf[1424] = f[657] && f[630] && f[633] && f[349]; // c8t948i94
	assign leaf[1425] = !f[571] && !f[595] && !f[569] && !f[513]; // c8t958i95
	assign leaf[1426] = !f[571] && !f[595] && !f[569] && f[513]; // c8t958i95
	assign leaf[1427] = !f[571] && !f[595] && f[569] && !f[494]; // c8t958i95
	assign leaf[1428] = !f[571] && !f[595] && f[569] && f[494]; // c8t958i95
	assign leaf[1429] = !f[571] && f[595] && !f[456] && !f[605]; // c8t958i95
	assign leaf[1430] = !f[571] && f[595] && !f[456] && f[605]; // c8t958i95
	assign leaf[1431] = !f[571] && f[595] && f[456] && !f[325]; // c8t958i95
	assign leaf[1432] = !f[571] && f[595] && f[456] && f[325]; // c8t958i95
	assign leaf[1433] = f[571] && !f[680] && !f[569] && !f[216]; // c8t958i95
	assign leaf[1434] = f[571] && !f[680] && !f[569] && f[216]; // c8t958i95
	assign leaf[1435] = f[571] && !f[680] && f[569] && !f[158]; // c8t958i95
	assign leaf[1436] = f[571] && !f[680] && f[569] && f[158]; // c8t958i95
	assign leaf[1437] = f[571] && f[680] && !f[683] && !f[541]; // c8t958i95
	assign leaf[1438] = f[571] && f[680] && !f[683] && f[541]; // c8t958i95
	assign leaf[1439] = f[571] && f[680] && f[683] && !f[569]; // c8t958i95
	assign leaf[1440] = f[571] && f[680] && f[683] && f[569]; // c8t958i95
	assign leaf[1441] = !f[442] && !f[258] && !f[526] && !f[601]; // c8t968i96
	assign leaf[1442] = !f[442] && !f[258] && !f[526] && f[601]; // c8t968i96
	assign leaf[1443] = !f[442] && !f[258] && f[526] && !f[484]; // c8t968i96
	assign leaf[1444] = !f[442] && !f[258] && f[526] && f[484]; // c8t968i96
	assign leaf[1445] = !f[442] && f[258] && !f[682] && !f[633]; // c8t968i96
	assign leaf[1446] = !f[442] && f[258] && !f[682] && f[633]; // c8t968i96
	assign leaf[1447] = !f[442] && f[258] && f[682]; // c8t968i96
	assign leaf[1448] = f[442] && !f[291] && !f[211]; // c8t968i96
	assign leaf[1449] = f[442] && !f[291] && f[211] && !f[598]; // c8t968i96
	assign leaf[1450] = f[442] && !f[291] && f[211] && f[598]; // c8t968i96
	assign leaf[1451] = f[442] && f[291] && !f[386]; // c8t968i96
	assign leaf[1452] = f[442] && f[291] && f[386]; // c8t968i96
	assign leaf[1453] = !f[211] && !f[636] && !f[154] && !f[569]; // c8t978i97
	assign leaf[1454] = !f[211] && !f[636] && !f[154] && f[569]; // c8t978i97
	assign leaf[1455] = !f[211] && !f[636] && f[154] && !f[322]; // c8t978i97
	assign leaf[1456] = !f[211] && !f[636] && f[154] && f[322]; // c8t978i97
	assign leaf[1457] = !f[211] && f[636] && !f[578] && !f[128]; // c8t978i97
	assign leaf[1458] = !f[211] && f[636] && !f[578] && f[128]; // c8t978i97
	assign leaf[1459] = !f[211] && f[636] && f[578] && !f[572]; // c8t978i97
	assign leaf[1460] = !f[211] && f[636] && f[578] && f[572]; // c8t978i97
	assign leaf[1461] = f[211] && !f[210] && !f[594] && !f[431]; // c8t978i97
	assign leaf[1462] = f[211] && !f[210] && !f[594] && f[431]; // c8t978i97
	assign leaf[1463] = f[211] && !f[210] && f[594] && !f[463]; // c8t978i97
	assign leaf[1464] = f[211] && !f[210] && f[594] && f[463]; // c8t978i97
	assign leaf[1465] = f[211] && f[210] && !f[263] && !f[273]; // c8t978i97
	assign leaf[1466] = f[211] && f[210] && !f[263] && f[273]; // c8t978i97
	assign leaf[1467] = f[211] && f[210] && f[263] && !f[204]; // c8t978i97
	assign leaf[1468] = f[211] && f[210] && f[263] && f[204]; // c8t978i97
	assign leaf[1469] = !f[458] && !f[512] && !f[488] && !f[517]; // c8t988i98
	assign leaf[1470] = !f[458] && !f[512] && !f[488] && f[517]; // c8t988i98
	assign leaf[1471] = !f[458] && !f[512] && f[488] && !f[517]; // c8t988i98
	assign leaf[1472] = !f[458] && !f[512] && f[488] && f[517]; // c8t988i98
	assign leaf[1473] = !f[458] && f[512] && !f[576] && !f[348]; // c8t988i98
	assign leaf[1474] = !f[458] && f[512] && !f[576] && f[348]; // c8t988i98
	assign leaf[1475] = !f[458] && f[512] && f[576] && !f[274]; // c8t988i98
	assign leaf[1476] = !f[458] && f[512] && f[576] && f[274]; // c8t988i98
	assign leaf[1477] = f[458] && !f[489] && !f[454] && !f[294]; // c8t988i98
	assign leaf[1478] = f[458] && !f[489] && !f[454] && f[294]; // c8t988i98
	assign leaf[1479] = f[458] && !f[489] && f[454] && !f[436]; // c8t988i98
	assign leaf[1480] = f[458] && !f[489] && f[454] && f[436]; // c8t988i98
	assign leaf[1481] = f[458] && f[489] && !f[373] && !f[596]; // c8t988i98
	assign leaf[1482] = f[458] && f[489] && !f[373] && f[596]; // c8t988i98
	assign leaf[1483] = f[458] && f[489] && f[373] && !f[521]; // c8t988i98
	assign leaf[1484] = f[458] && f[489] && f[373] && f[521]; // c8t988i98
	assign leaf[1485] = !f[303] && !f[594] && !f[650] && !f[271]; // c8t998i99
	assign leaf[1486] = !f[303] && !f[594] && !f[650] && f[271]; // c8t998i99
	assign leaf[1487] = !f[303] && !f[594] && f[650] && !f[601]; // c8t998i99
	assign leaf[1488] = !f[303] && !f[594] && f[650] && f[601]; // c8t998i99
	assign leaf[1489] = !f[303] && f[594] && !f[463] && !f[465]; // c8t998i99
	assign leaf[1490] = !f[303] && f[594] && !f[463] && f[465]; // c8t998i99
	assign leaf[1491] = !f[303] && f[594] && f[463] && !f[487]; // c8t998i99
	assign leaf[1492] = !f[303] && f[594] && f[463] && f[487]; // c8t998i99
	assign leaf[1493] = f[303] && !f[649] && !f[682] && !f[207]; // c8t998i99
	assign leaf[1494] = f[303] && !f[649] && !f[682] && f[207]; // c8t998i99
	assign leaf[1495] = f[303] && !f[649] && f[682] && !f[595]; // c8t998i99
	assign leaf[1496] = f[303] && !f[649] && f[682] && f[595]; // c8t998i99
	assign leaf[1497] = f[303] && f[649]; // c8t998i99
endmodule

module decision_tree_leaves_9(input logic [0:783] f, output logic [0:1347] leaf);
	assign leaf[0] = !f[717] && !f[713] && !f[715] && !f[711]; // c9t9i0
	assign leaf[1] = !f[717] && !f[713] && !f[715] && f[711]; // c9t9i0
	assign leaf[2] = !f[717] && !f[713] && f[715] && !f[210]; // c9t9i0
	assign leaf[3] = !f[717] && !f[713] && f[715] && f[210]; // c9t9i0
	assign leaf[4] = !f[717] && f[713] && !f[430] && !f[375]; // c9t9i0
	assign leaf[5] = !f[717] && f[713] && !f[430] && f[375]; // c9t9i0
	assign leaf[6] = !f[717] && f[713] && f[430] && !f[211]; // c9t9i0
	assign leaf[7] = !f[717] && f[713] && f[430] && f[211]; // c9t9i0
	assign leaf[8] = f[717] && !f[210] && !f[208] && !f[459]; // c9t9i0
	assign leaf[9] = f[717] && !f[210] && !f[208] && f[459]; // c9t9i0
	assign leaf[10] = f[717] && !f[210] && f[208] && !f[378]; // c9t9i0
	assign leaf[11] = f[717] && !f[210] && f[208] && f[378]; // c9t9i0
	assign leaf[12] = f[717] && f[210] && !f[231] && !f[685]; // c9t9i0
	assign leaf[13] = f[717] && f[210] && !f[231] && f[685]; // c9t9i0
	assign leaf[14] = f[717] && f[210] && f[231] && !f[398]; // c9t9i0
	assign leaf[15] = f[717] && f[210] && f[231] && f[398]; // c9t9i0
	assign leaf[16] = !f[156] && !f[211] && !f[720] && !f[239]; // c9t19i1
	assign leaf[17] = !f[156] && !f[211] && !f[720] && f[239]; // c9t19i1
	assign leaf[18] = !f[156] && !f[211] && f[720] && !f[209]; // c9t19i1
	assign leaf[19] = !f[156] && !f[211] && f[720] && f[209]; // c9t19i1
	assign leaf[20] = !f[156] && f[211] && !f[409] && !f[408]; // c9t19i1
	assign leaf[21] = !f[156] && f[211] && !f[409] && f[408]; // c9t19i1
	assign leaf[22] = !f[156] && f[211] && f[409] && !f[345]; // c9t19i1
	assign leaf[23] = !f[156] && f[211] && f[409] && f[345]; // c9t19i1
	assign leaf[24] = f[156] && !f[128] && !f[409] && !f[439]; // c9t19i1
	assign leaf[25] = f[156] && !f[128] && !f[409] && f[439]; // c9t19i1
	assign leaf[26] = f[156] && !f[128] && f[409] && !f[626]; // c9t19i1
	assign leaf[27] = f[156] && !f[128] && f[409] && f[626]; // c9t19i1
	assign leaf[28] = f[156] && f[128] && !f[368]; // c9t19i1
	assign leaf[29] = f[156] && f[128] && f[368]; // c9t19i1
	assign leaf[30] = !f[597] && !f[381] && !f[721] && !f[383]; // c9t29i2
	assign leaf[31] = !f[597] && !f[381] && !f[721] && f[383]; // c9t29i2
	assign leaf[32] = !f[597] && !f[381] && f[721] && !f[488]; // c9t29i2
	assign leaf[33] = !f[597] && !f[381] && f[721] && f[488]; // c9t29i2
	assign leaf[34] = !f[597] && f[381] && !f[211] && !f[238]; // c9t29i2
	assign leaf[35] = !f[597] && f[381] && !f[211] && f[238]; // c9t29i2
	assign leaf[36] = !f[597] && f[381] && f[211] && !f[205]; // c9t29i2
	assign leaf[37] = !f[597] && f[381] && f[211] && f[205]; // c9t29i2
	assign leaf[38] = f[597] && !f[707] && !f[706] && !f[708]; // c9t29i2
	assign leaf[39] = f[597] && !f[707] && !f[706] && f[708]; // c9t29i2
	assign leaf[40] = f[597] && !f[707] && f[706]; // c9t29i2
	assign leaf[41] = f[597] && f[707] && !f[376] && !f[429]; // c9t29i2
	assign leaf[42] = f[597] && f[707] && !f[376] && f[429]; // c9t29i2
	assign leaf[43] = f[597] && f[707] && f[376] && !f[219]; // c9t29i2
	assign leaf[44] = f[597] && f[707] && f[376] && f[219]; // c9t29i2
	assign leaf[45] = !f[569] && !f[381] && !f[342] && !f[290]; // c9t39i3
	assign leaf[46] = !f[569] && !f[381] && !f[342] && f[290]; // c9t39i3
	assign leaf[47] = !f[569] && !f[381] && f[342] && !f[209]; // c9t39i3
	assign leaf[48] = !f[569] && !f[381] && f[342] && f[209]; // c9t39i3
	assign leaf[49] = !f[569] && f[381] && !f[211] && !f[239]; // c9t39i3
	assign leaf[50] = !f[569] && f[381] && !f[211] && f[239]; // c9t39i3
	assign leaf[51] = !f[569] && f[381] && f[211] && !f[155]; // c9t39i3
	assign leaf[52] = !f[569] && f[381] && f[211] && f[155]; // c9t39i3
	assign leaf[53] = f[569] && !f[692] && !f[706] && !f[707]; // c9t39i3
	assign leaf[54] = f[569] && !f[692] && !f[706] && f[707]; // c9t39i3
	assign leaf[55] = f[569] && !f[692] && f[706] && !f[377]; // c9t39i3
	assign leaf[56] = f[569] && !f[692] && f[706] && f[377]; // c9t39i3
	assign leaf[57] = f[569] && f[692] && !f[482] && !f[511]; // c9t39i3
	assign leaf[58] = f[569] && f[692] && !f[482] && f[511]; // c9t39i3
	assign leaf[59] = f[569] && f[692] && f[482]; // c9t39i3
	assign leaf[60] = !f[598] && !f[372] && !f[398] && !f[346]; // c9t49i4
	assign leaf[61] = !f[598] && !f[372] && !f[398] && f[346]; // c9t49i4
	assign leaf[62] = !f[598] && !f[372] && f[398] && !f[209]; // c9t49i4
	assign leaf[63] = !f[598] && !f[372] && f[398] && f[209]; // c9t49i4
	assign leaf[64] = !f[598] && f[372] && !f[210] && !f[238]; // c9t49i4
	assign leaf[65] = !f[598] && f[372] && !f[210] && f[238]; // c9t49i4
	assign leaf[66] = !f[598] && f[372] && f[210] && !f[347]; // c9t49i4
	assign leaf[67] = !f[598] && f[372] && f[210] && f[347]; // c9t49i4
	assign leaf[68] = f[598] && !f[708] && !f[706] && !f[709]; // c9t49i4
	assign leaf[69] = f[598] && !f[708] && !f[706] && f[709]; // c9t49i4
	assign leaf[70] = f[598] && !f[708] && f[706] && !f[406]; // c9t49i4
	assign leaf[71] = f[598] && !f[708] && f[706] && f[406]; // c9t49i4
	assign leaf[72] = f[598] && f[708] && !f[405] && !f[350]; // c9t49i4
	assign leaf[73] = f[598] && f[708] && !f[405] && f[350]; // c9t49i4
	assign leaf[74] = f[598] && f[708] && f[405] && !f[233]; // c9t49i4
	assign leaf[75] = f[598] && f[708] && f[405] && f[233]; // c9t49i4
	assign leaf[76] = !f[570] && !f[624] && !f[212] && !f[692]; // c9t59i5
	assign leaf[77] = !f[570] && !f[624] && !f[212] && f[692]; // c9t59i5
	assign leaf[78] = !f[570] && !f[624] && f[212] && !f[205]; // c9t59i5
	assign leaf[79] = !f[570] && !f[624] && f[212] && f[205]; // c9t59i5
	assign leaf[80] = !f[570] && f[624] && !f[706] && !f[238]; // c9t59i5
	assign leaf[81] = !f[570] && f[624] && !f[706] && f[238]; // c9t59i5
	assign leaf[82] = !f[570] && f[624] && f[706]; // c9t59i5
	assign leaf[83] = f[570] && !f[680] && !f[719] && !f[340]; // c9t59i5
	assign leaf[84] = f[570] && !f[680] && !f[719] && f[340]; // c9t59i5
	assign leaf[85] = f[570] && !f[680] && f[719] && !f[573]; // c9t59i5
	assign leaf[86] = f[570] && !f[680] && f[719] && f[573]; // c9t59i5
	assign leaf[87] = f[570] && f[680] && !f[374] && !f[348]; // c9t59i5
	assign leaf[88] = f[570] && f[680] && !f[374] && f[348]; // c9t59i5
	assign leaf[89] = f[570] && f[680] && f[374] && !f[214]; // c9t59i5
	assign leaf[90] = f[570] && f[680] && f[374] && f[214]; // c9t59i5
	assign leaf[91] = !f[569] && !f[354] && !f[157] && !f[290]; // c9t69i6
	assign leaf[92] = !f[569] && !f[354] && !f[157] && f[290]; // c9t69i6
	assign leaf[93] = !f[569] && !f[354] && f[157] && !f[384]; // c9t69i6
	assign leaf[94] = !f[569] && !f[354] && f[157] && f[384]; // c9t69i6
	assign leaf[95] = !f[569] && f[354] && !f[406] && !f[487]; // c9t69i6
	assign leaf[96] = !f[569] && f[354] && !f[406] && f[487]; // c9t69i6
	assign leaf[97] = !f[569] && f[354] && f[406] && !f[623]; // c9t69i6
	assign leaf[98] = !f[569] && f[354] && f[406] && f[623]; // c9t69i6
	assign leaf[99] = f[569] && !f[368] && !f[706] && !f[689]; // c9t69i6
	assign leaf[100] = f[569] && !f[368] && !f[706] && f[689]; // c9t69i6
	assign leaf[101] = f[569] && !f[368] && f[706] && !f[376]; // c9t69i6
	assign leaf[102] = f[569] && !f[368] && f[706] && f[376]; // c9t69i6
	assign leaf[103] = f[569] && f[368] && !f[355]; // c9t69i6
	assign leaf[104] = f[569] && f[368] && f[355] && !f[340]; // c9t69i6
	assign leaf[105] = f[569] && f[368] && f[355] && f[340]; // c9t69i6
	assign leaf[106] = !f[570] && !f[624] && !f[212] && !f[719]; // c9t79i7
	assign leaf[107] = !f[570] && !f[624] && !f[212] && f[719]; // c9t79i7
	assign leaf[108] = !f[570] && !f[624] && f[212] && !f[204]; // c9t79i7
	assign leaf[109] = !f[570] && !f[624] && f[212] && f[204]; // c9t79i7
	assign leaf[110] = !f[570] && f[624] && !f[384] && !f[324]; // c9t79i7
	assign leaf[111] = !f[570] && f[624] && !f[384] && f[324]; // c9t79i7
	assign leaf[112] = !f[570] && f[624] && f[384] && !f[680]; // c9t79i7
	assign leaf[113] = !f[570] && f[624] && f[384] && f[680]; // c9t79i7
	assign leaf[114] = f[570] && !f[680] && !f[720] && !f[599]; // c9t79i7
	assign leaf[115] = f[570] && !f[680] && !f[720] && f[599]; // c9t79i7
	assign leaf[116] = f[570] && !f[680] && f[720]; // c9t79i7
	assign leaf[117] = f[570] && f[680] && !f[207] && !f[213]; // c9t79i7
	assign leaf[118] = f[570] && f[680] && !f[207] && f[213]; // c9t79i7
	assign leaf[119] = f[570] && f[680] && f[207] && !f[377]; // c9t79i7
	assign leaf[120] = f[570] && f[680] && f[207] && f[377]; // c9t79i7
	assign leaf[121] = !f[157] && !f[571] && !f[203] && !f[189]; // c9t89i8
	assign leaf[122] = !f[157] && !f[571] && !f[203] && f[189]; // c9t89i8
	assign leaf[123] = !f[157] && !f[571] && f[203] && !f[342]; // c9t89i8
	assign leaf[124] = !f[157] && !f[571] && f[203] && f[342]; // c9t89i8
	assign leaf[125] = !f[157] && f[571] && !f[709] && !f[679]; // c9t89i8
	assign leaf[126] = !f[157] && f[571] && !f[709] && f[679]; // c9t89i8
	assign leaf[127] = !f[157] && f[571] && f[709] && !f[185]; // c9t89i8
	assign leaf[128] = !f[157] && f[571] && f[709] && f[185]; // c9t89i8
	assign leaf[129] = f[157] && !f[372] && !f[397] && !f[291]; // c9t89i8
	assign leaf[130] = f[157] && !f[372] && !f[397] && f[291]; // c9t89i8
	assign leaf[131] = f[157] && !f[372] && f[397] && !f[552]; // c9t89i8
	assign leaf[132] = f[157] && !f[372] && f[397] && f[552]; // c9t89i8
	assign leaf[133] = f[157] && f[372] && !f[235] && !f[236]; // c9t89i8
	assign leaf[134] = f[157] && f[372] && !f[235] && f[236]; // c9t89i8
	assign leaf[135] = f[157] && f[372] && f[235] && !f[552]; // c9t89i8
	assign leaf[136] = f[157] && f[372] && f[235] && f[552]; // c9t89i8
	assign leaf[137] = !f[154] && !f[596] && !f[210] && !f[266]; // c9t99i9
	assign leaf[138] = !f[154] && !f[596] && !f[210] && f[266]; // c9t99i9
	assign leaf[139] = !f[154] && !f[596] && f[210] && !f[206]; // c9t99i9
	assign leaf[140] = !f[154] && !f[596] && f[210] && f[206]; // c9t99i9
	assign leaf[141] = !f[154] && f[596] && !f[706] && !f[665]; // c9t99i9
	assign leaf[142] = !f[154] && f[596] && !f[706] && f[665]; // c9t99i9
	assign leaf[143] = !f[154] && f[596] && f[706] && !f[375]; // c9t99i9
	assign leaf[144] = !f[154] && f[596] && f[706] && f[375]; // c9t99i9
	assign leaf[145] = f[154] && !f[316] && !f[290] && !f[342]; // c9t99i9
	assign leaf[146] = f[154] && !f[316] && !f[290] && f[342]; // c9t99i9
	assign leaf[147] = f[154] && !f[316] && f[290] && !f[571]; // c9t99i9
	assign leaf[148] = f[154] && !f[316] && f[290] && f[571]; // c9t99i9
	assign leaf[149] = f[154] && f[316] && !f[600] && !f[354]; // c9t99i9
	assign leaf[150] = f[154] && f[316] && !f[600] && f[354]; // c9t99i9
	assign leaf[151] = f[154] && f[316] && f[600] && !f[544]; // c9t99i9
	assign leaf[152] = f[154] && f[316] && f[600] && f[544]; // c9t99i9
	assign leaf[153] = !f[568] && !f[720] && !f[177] && !f[294]; // c9t109i10
	assign leaf[154] = !f[568] && !f[720] && !f[177] && f[294]; // c9t109i10
	assign leaf[155] = !f[568] && !f[720] && f[177] && !f[287]; // c9t109i10
	assign leaf[156] = !f[568] && !f[720] && f[177] && f[287]; // c9t109i10
	assign leaf[157] = !f[568] && f[720] && !f[717] && !f[202]; // c9t109i10
	assign leaf[158] = !f[568] && f[720] && !f[717] && f[202]; // c9t109i10
	assign leaf[159] = !f[568] && f[720] && f[717] && !f[429]; // c9t109i10
	assign leaf[160] = !f[568] && f[720] && f[717] && f[429]; // c9t109i10
	assign leaf[161] = f[568] && !f[341] && !f[689] && !f[676]; // c9t109i10
	assign leaf[162] = f[568] && !f[341] && !f[689] && f[676]; // c9t109i10
	assign leaf[163] = f[568] && !f[341] && f[689] && !f[625]; // c9t109i10
	assign leaf[164] = f[568] && !f[341] && f[689] && f[625]; // c9t109i10
	assign leaf[165] = f[568] && f[341] && !f[543] && !f[573]; // c9t109i10
	assign leaf[166] = f[568] && f[341] && !f[543] && f[573]; // c9t109i10
	assign leaf[167] = f[568] && f[341] && f[543] && !f[576]; // c9t109i10
	assign leaf[168] = f[568] && f[341] && f[543] && f[576]; // c9t109i10
	assign leaf[169] = !f[158] && !f[126] && !f[218] && !f[400]; // c9t119i11
	assign leaf[170] = !f[158] && !f[126] && !f[218] && f[400]; // c9t119i11
	assign leaf[171] = !f[158] && !f[126] && f[218] && !f[214]; // c9t119i11
	assign leaf[172] = !f[158] && !f[126] && f[218] && f[214]; // c9t119i11
	assign leaf[173] = !f[158] && f[126] && !f[626]; // c9t119i11
	assign leaf[174] = !f[158] && f[126] && f[626] && !f[261]; // c9t119i11
	assign leaf[175] = !f[158] && f[126] && f[626] && f[261]; // c9t119i11
	assign leaf[176] = f[158] && !f[329] && !f[518] && !f[356]; // c9t119i11
	assign leaf[177] = f[158] && !f[329] && !f[518] && f[356]; // c9t119i11
	assign leaf[178] = f[158] && !f[329] && f[518] && !f[241]; // c9t119i11
	assign leaf[179] = f[158] && !f[329] && f[518] && f[241]; // c9t119i11
	assign leaf[180] = f[158] && f[329] && !f[372] && !f[371]; // c9t119i11
	assign leaf[181] = f[158] && f[329] && !f[372] && f[371]; // c9t119i11
	assign leaf[182] = f[158] && f[329] && f[372] && !f[411]; // c9t119i11
	assign leaf[183] = f[158] && f[329] && f[372] && f[411]; // c9t119i11
	assign leaf[184] = !f[719] && !f[578] && !f[318] && !f[316]; // c9t129i12
	assign leaf[185] = !f[719] && !f[578] && !f[318] && f[316]; // c9t129i12
	assign leaf[186] = !f[719] && !f[578] && f[318] && !f[468]; // c9t129i12
	assign leaf[187] = !f[719] && !f[578] && f[318] && f[468]; // c9t129i12
	assign leaf[188] = !f[719] && f[578] && !f[399] && !f[718]; // c9t129i12
	assign leaf[189] = !f[719] && f[578] && !f[399] && f[718]; // c9t129i12
	assign leaf[190] = !f[719] && f[578] && f[399] && !f[346]; // c9t129i12
	assign leaf[191] = !f[719] && f[578] && f[399] && f[346]; // c9t129i12
	assign leaf[192] = f[719] && !f[717] && !f[201] && !f[319]; // c9t129i12
	assign leaf[193] = f[719] && !f[717] && !f[201] && f[319]; // c9t129i12
	assign leaf[194] = f[719] && !f[717] && f[201] && !f[459]; // c9t129i12
	assign leaf[195] = f[719] && !f[717] && f[201] && f[459]; // c9t129i12
	assign leaf[196] = f[719] && f[717] && !f[431] && !f[458]; // c9t129i12
	assign leaf[197] = f[719] && f[717] && !f[431] && f[458]; // c9t129i12
	assign leaf[198] = f[719] && f[717] && f[431] && !f[633]; // c9t129i12
	assign leaf[199] = f[719] && f[717] && f[431] && f[633]; // c9t129i12
	assign leaf[200] = !f[159] && !f[632] && !f[212] && !f[572]; // c9t139i13
	assign leaf[201] = !f[159] && !f[632] && !f[212] && f[572]; // c9t139i13
	assign leaf[202] = !f[159] && !f[632] && f[212] && !f[291]; // c9t139i13
	assign leaf[203] = !f[159] && !f[632] && f[212] && f[291]; // c9t139i13
	assign leaf[204] = !f[159] && f[632] && !f[601] && !f[683]; // c9t139i13
	assign leaf[205] = !f[159] && f[632] && !f[601] && f[683]; // c9t139i13
	assign leaf[206] = !f[159] && f[632] && f[601] && !f[517]; // c9t139i13
	assign leaf[207] = !f[159] && f[632] && f[601] && f[517]; // c9t139i13
	assign leaf[208] = f[159] && !f[355] && !f[657] && !f[688]; // c9t139i13
	assign leaf[209] = f[159] && !f[355] && !f[657] && f[688]; // c9t139i13
	assign leaf[210] = f[159] && !f[355] && f[657]; // c9t139i13
	assign leaf[211] = f[159] && f[355] && !f[290] && !f[682]; // c9t139i13
	assign leaf[212] = f[159] && f[355] && !f[290] && f[682]; // c9t139i13
	assign leaf[213] = f[159] && f[355] && f[290] && !f[493]; // c9t139i13
	assign leaf[214] = f[159] && f[355] && f[290] && f[493]; // c9t139i13
	assign leaf[215] = !f[469] && !f[436] && !f[438] && !f[468]; // c9t149i14
	assign leaf[216] = !f[469] && !f[436] && !f[438] && f[468]; // c9t149i14
	assign leaf[217] = !f[469] && !f[436] && f[438] && !f[320]; // c9t149i14
	assign leaf[218] = !f[469] && !f[436] && f[438] && f[320]; // c9t149i14
	assign leaf[219] = !f[469] && f[436] && !f[567] && !f[233]; // c9t149i14
	assign leaf[220] = !f[469] && f[436] && !f[567] && f[233]; // c9t149i14
	assign leaf[221] = !f[469] && f[436] && f[567] && !f[398]; // c9t149i14
	assign leaf[222] = !f[469] && f[436] && f[567] && f[398]; // c9t149i14
	assign leaf[223] = f[469] && !f[369] && !f[694] && !f[385]; // c9t149i14
	assign leaf[224] = f[469] && !f[369] && !f[694] && f[385]; // c9t149i14
	assign leaf[225] = f[469] && !f[369] && f[694]; // c9t149i14
	assign leaf[226] = f[469] && f[369] && !f[385] && !f[667]; // c9t149i14
	assign leaf[227] = f[469] && f[369] && !f[385] && f[667]; // c9t149i14
	assign leaf[228] = f[469] && f[369] && f[385] && !f[229]; // c9t149i14
	assign leaf[229] = f[469] && f[369] && f[385] && f[229]; // c9t149i14
	assign leaf[230] = !f[128] && !f[443] && !f[189] && !f[355]; // c9t159i15
	assign leaf[231] = !f[128] && !f[443] && !f[189] && f[355]; // c9t159i15
	assign leaf[232] = !f[128] && !f[443] && f[189] && !f[383]; // c9t159i15
	assign leaf[233] = !f[128] && !f[443] && f[189] && f[383]; // c9t159i15
	assign leaf[234] = !f[128] && f[443] && !f[639] && !f[368]; // c9t159i15
	assign leaf[235] = !f[128] && f[443] && !f[639] && f[368]; // c9t159i15
	assign leaf[236] = !f[128] && f[443] && f[639]; // c9t159i15
	assign leaf[237] = f[128] && !f[275] && !f[659] && !f[358]; // c9t159i15
	assign leaf[238] = f[128] && !f[275] && !f[659] && f[358]; // c9t159i15
	assign leaf[239] = f[128] && !f[275] && f[659] && !f[432]; // c9t159i15
	assign leaf[240] = f[128] && !f[275] && f[659] && f[432]; // c9t159i15
	assign leaf[241] = f[128] && f[275]; // c9t159i15
	assign leaf[242] = !f[160] && !f[176] && !f[126] && !f[219]; // c9t169i16
	assign leaf[243] = !f[160] && !f[176] && !f[126] && f[219]; // c9t169i16
	assign leaf[244] = !f[160] && !f[176] && f[126] && !f[462]; // c9t169i16
	assign leaf[245] = !f[160] && !f[176] && f[126] && f[462]; // c9t169i16
	assign leaf[246] = !f[160] && f[176] && !f[694] && !f[342]; // c9t169i16
	assign leaf[247] = !f[160] && f[176] && !f[694] && f[342]; // c9t169i16
	assign leaf[248] = !f[160] && f[176] && f[694] && !f[440]; // c9t169i16
	assign leaf[249] = !f[160] && f[176] && f[694] && f[440]; // c9t169i16
	assign leaf[250] = f[160] && !f[427] && !f[572] && !f[509]; // c9t169i16
	assign leaf[251] = f[160] && !f[427] && !f[572] && f[509]; // c9t169i16
	assign leaf[252] = f[160] && !f[427] && f[572] && !f[318]; // c9t169i16
	assign leaf[253] = f[160] && !f[427] && f[572] && f[318]; // c9t169i16
	assign leaf[254] = f[160] && f[427] && !f[264]; // c9t169i16
	assign leaf[255] = f[160] && f[427] && f[264] && !f[595]; // c9t169i16
	assign leaf[256] = f[160] && f[427] && f[264] && f[595]; // c9t169i16
	assign leaf[257] = !f[694] && !f[742] && !f[719] && !f[380]; // c9t179i17
	assign leaf[258] = !f[694] && !f[742] && !f[719] && f[380]; // c9t179i17
	assign leaf[259] = !f[694] && !f[742] && f[719] && !f[659]; // c9t179i17
	assign leaf[260] = !f[694] && !f[742] && f[719] && f[659]; // c9t179i17
	assign leaf[261] = !f[694] && f[742] && !f[259] && !f[350]; // c9t179i17
	assign leaf[262] = !f[694] && f[742] && !f[259] && f[350]; // c9t179i17
	assign leaf[263] = !f[694] && f[742] && f[259] && !f[329]; // c9t179i17
	assign leaf[264] = !f[694] && f[742] && f[259] && f[329]; // c9t179i17
	assign leaf[265] = f[694] && !f[439] && !f[465]; // c9t179i17
	assign leaf[266] = f[694] && !f[439] && f[465] && !f[314]; // c9t179i17
	assign leaf[267] = f[694] && !f[439] && f[465] && f[314]; // c9t179i17
	assign leaf[268] = f[694] && f[439] && !f[174] && !f[216]; // c9t179i17
	assign leaf[269] = f[694] && f[439] && !f[174] && f[216]; // c9t179i17
	assign leaf[270] = f[694] && f[439] && f[174]; // c9t179i17
	assign leaf[271] = !f[159] && !f[203] && !f[742] && !f[692]; // c9t189i18
	assign leaf[272] = !f[159] && !f[203] && !f[742] && f[692]; // c9t189i18
	assign leaf[273] = !f[159] && !f[203] && f[742] && !f[232]; // c9t189i18
	assign leaf[274] = !f[159] && !f[203] && f[742] && f[232]; // c9t189i18
	assign leaf[275] = !f[159] && f[203] && !f[314] && !f[397]; // c9t189i18
	assign leaf[276] = !f[159] && f[203] && !f[314] && f[397]; // c9t189i18
	assign leaf[277] = !f[159] && f[203] && f[314] && !f[206]; // c9t189i18
	assign leaf[278] = !f[159] && f[203] && f[314] && f[206]; // c9t189i18
	assign leaf[279] = f[159] && !f[357] && !f[346] && !f[689]; // c9t189i18
	assign leaf[280] = f[159] && !f[357] && !f[346] && f[689]; // c9t189i18
	assign leaf[281] = f[159] && !f[357] && f[346] && !f[549]; // c9t189i18
	assign leaf[282] = f[159] && !f[357] && f[346] && f[549]; // c9t189i18
	assign leaf[283] = f[159] && f[357] && !f[439]; // c9t189i18
	assign leaf[284] = f[159] && f[357] && f[439] && !f[262]; // c9t189i18
	assign leaf[285] = f[159] && f[357] && f[439] && f[262]; // c9t189i18
	assign leaf[286] = !f[567] && !f[659] && !f[212] && !f[545]; // c9t199i19
	assign leaf[287] = !f[567] && !f[659] && !f[212] && f[545]; // c9t199i19
	assign leaf[288] = !f[567] && !f[659] && f[212] && !f[327]; // c9t199i19
	assign leaf[289] = !f[567] && !f[659] && f[212] && f[327]; // c9t199i19
	assign leaf[290] = !f[567] && f[659] && !f[545] && !f[742]; // c9t199i19
	assign leaf[291] = !f[567] && f[659] && !f[545] && f[742]; // c9t199i19
	assign leaf[292] = !f[567] && f[659] && f[545] && !f[485]; // c9t199i19
	assign leaf[293] = !f[567] && f[659] && f[545] && f[485]; // c9t199i19
	assign leaf[294] = f[567] && !f[369] && !f[485] && !f[566]; // c9t199i19
	assign leaf[295] = f[567] && !f[369] && !f[485] && f[566]; // c9t199i19
	assign leaf[296] = f[567] && !f[369] && f[485] && !f[399]; // c9t199i19
	assign leaf[297] = f[567] && !f[369] && f[485] && f[399]; // c9t199i19
	assign leaf[298] = f[567] && f[369] && !f[471] && !f[466]; // c9t199i19
	assign leaf[299] = f[567] && f[369] && !f[471] && f[466]; // c9t199i19
	assign leaf[300] = f[567] && f[369] && f[471]; // c9t199i19
	assign leaf[301] = !f[599] && !f[229] && !f[653] && !f[443]; // c9t209i20
	assign leaf[302] = !f[599] && !f[229] && !f[653] && f[443]; // c9t209i20
	assign leaf[303] = !f[599] && !f[229] && f[653] && !f[155]; // c9t209i20
	assign leaf[304] = !f[599] && !f[229] && f[653] && f[155]; // c9t209i20
	assign leaf[305] = !f[599] && f[229] && !f[177] && !f[205]; // c9t209i20
	assign leaf[306] = !f[599] && f[229] && !f[177] && f[205]; // c9t209i20
	assign leaf[307] = !f[599] && f[229] && f[177] && !f[183]; // c9t209i20
	assign leaf[308] = !f[599] && f[229] && f[177] && f[183]; // c9t209i20
	assign leaf[309] = f[599] && !f[709] && !f[680] && !f[543]; // c9t209i20
	assign leaf[310] = f[599] && !f[709] && !f[680] && f[543]; // c9t209i20
	assign leaf[311] = f[599] && !f[709] && f[680] && !f[207]; // c9t209i20
	assign leaf[312] = f[599] && !f[709] && f[680] && f[207]; // c9t209i20
	assign leaf[313] = f[599] && f[709] && !f[235] && !f[214]; // c9t209i20
	assign leaf[314] = f[599] && f[709] && !f[235] && f[214]; // c9t209i20
	assign leaf[315] = f[599] && f[709] && f[235] && !f[378]; // c9t209i20
	assign leaf[316] = f[599] && f[709] && f[235] && f[378]; // c9t209i20
	assign leaf[317] = !f[150] && !f[129] && !f[191] && !f[355]; // c9t219i21
	assign leaf[318] = !f[150] && !f[129] && !f[191] && f[355]; // c9t219i21
	assign leaf[319] = !f[150] && !f[129] && f[191] && !f[187]; // c9t219i21
	assign leaf[320] = !f[150] && !f[129] && f[191] && f[187]; // c9t219i21
	assign leaf[321] = !f[150] && f[129] && !f[126] && !f[609]; // c9t219i21
	assign leaf[322] = !f[150] && f[129] && !f[126] && f[609]; // c9t219i21
	assign leaf[323] = !f[150] && f[129] && f[126] && !f[289]; // c9t219i21
	assign leaf[324] = !f[150] && f[129] && f[126] && f[289]; // c9t219i21
	assign leaf[325] = f[150] && !f[259] && !f[685] && !f[686]; // c9t219i21
	assign leaf[326] = f[150] && !f[259] && !f[685] && f[686]; // c9t219i21
	assign leaf[327] = f[150] && !f[259] && f[685] && !f[411]; // c9t219i21
	assign leaf[328] = f[150] && !f[259] && f[685] && f[411]; // c9t219i21
	assign leaf[329] = f[150] && f[259] && !f[522] && !f[267]; // c9t219i21
	assign leaf[330] = f[150] && f[259] && !f[522] && f[267]; // c9t219i21
	assign leaf[331] = f[150] && f[259] && f[522] && !f[464]; // c9t219i21
	assign leaf[332] = f[150] && f[259] && f[522] && f[464]; // c9t219i21
	assign leaf[333] = !f[469] && !f[353] && !f[405] && !f[455]; // c9t229i22
	assign leaf[334] = !f[469] && !f[353] && !f[405] && f[455]; // c9t229i22
	assign leaf[335] = !f[469] && !f[353] && f[405] && !f[660]; // c9t229i22
	assign leaf[336] = !f[469] && !f[353] && f[405] && f[660]; // c9t229i22
	assign leaf[337] = !f[469] && f[353] && !f[378] && !f[350]; // c9t229i22
	assign leaf[338] = !f[469] && f[353] && !f[378] && f[350]; // c9t229i22
	assign leaf[339] = !f[469] && f[353] && f[378] && !f[461]; // c9t229i22
	assign leaf[340] = !f[469] && f[353] && f[378] && f[461]; // c9t229i22
	assign leaf[341] = f[469] && !f[385] && !f[667] && !f[720]; // c9t229i22
	assign leaf[342] = f[469] && !f[385] && !f[667] && f[720]; // c9t229i22
	assign leaf[343] = f[469] && !f[385] && f[667]; // c9t229i22
	assign leaf[344] = f[469] && f[385] && !f[313] && !f[470]; // c9t229i22
	assign leaf[345] = f[469] && f[385] && !f[313] && f[470]; // c9t229i22
	assign leaf[346] = f[469] && f[385] && f[313] && !f[182]; // c9t229i22
	assign leaf[347] = f[469] && f[385] && f[313] && f[182]; // c9t229i22
	assign leaf[348] = !f[571] && !f[188] && !f[218] && !f[378]; // c9t239i23
	assign leaf[349] = !f[571] && !f[188] && !f[218] && f[378]; // c9t239i23
	assign leaf[350] = !f[571] && !f[188] && f[218] && !f[211]; // c9t239i23
	assign leaf[351] = !f[571] && !f[188] && f[218] && f[211]; // c9t239i23
	assign leaf[352] = !f[571] && f[188] && !f[383] && !f[545]; // c9t239i23
	assign leaf[353] = !f[571] && f[188] && !f[383] && f[545]; // c9t239i23
	assign leaf[354] = !f[571] && f[188] && f[383] && !f[574]; // c9t239i23
	assign leaf[355] = !f[571] && f[188] && f[383] && f[574]; // c9t239i23
	assign leaf[356] = f[571] && !f[213] && !f[425] && !f[574]; // c9t239i23
	assign leaf[357] = f[571] && !f[213] && !f[425] && f[574]; // c9t239i23
	assign leaf[358] = f[571] && !f[213] && f[425] && !f[240]; // c9t239i23
	assign leaf[359] = f[571] && !f[213] && f[425] && f[240]; // c9t239i23
	assign leaf[360] = f[571] && f[213] && !f[657] && !f[319]; // c9t239i23
	assign leaf[361] = f[571] && f[213] && !f[657] && f[319]; // c9t239i23
	assign leaf[362] = f[571] && f[213] && f[657] && !f[488]; // c9t239i23
	assign leaf[363] = f[571] && f[213] && f[657] && f[488]; // c9t239i23
	assign leaf[364] = !f[571] && !f[443] && !f[569] && !f[176]; // c9t249i24
	assign leaf[365] = !f[571] && !f[443] && !f[569] && f[176]; // c9t249i24
	assign leaf[366] = !f[571] && !f[443] && f[569] && !f[486]; // c9t249i24
	assign leaf[367] = !f[571] && !f[443] && f[569] && f[486]; // c9t249i24
	assign leaf[368] = !f[571] && f[443] && !f[368] && !f[683]; // c9t249i24
	assign leaf[369] = !f[571] && f[443] && !f[368] && f[683]; // c9t249i24
	assign leaf[370] = !f[571] && f[443] && f[368]; // c9t249i24
	assign leaf[371] = f[571] && !f[680] && !f[488] && !f[213]; // c9t249i24
	assign leaf[372] = f[571] && !f[680] && !f[488] && f[213]; // c9t249i24
	assign leaf[373] = f[571] && !f[680] && f[488] && !f[678]; // c9t249i24
	assign leaf[374] = f[571] && !f[680] && f[488] && f[678]; // c9t249i24
	assign leaf[375] = f[571] && f[680] && !f[207] && !f[215]; // c9t249i24
	assign leaf[376] = f[571] && f[680] && !f[207] && f[215]; // c9t249i24
	assign leaf[377] = f[571] && f[680] && f[207] && !f[345]; // c9t249i24
	assign leaf[378] = f[571] && f[680] && f[207] && f[345]; // c9t249i24
	assign leaf[379] = !f[544] && !f[380] && !f[488] && !f[324]; // c9t259i25
	assign leaf[380] = !f[544] && !f[380] && !f[488] && f[324]; // c9t259i25
	assign leaf[381] = !f[544] && !f[380] && f[488] && !f[348]; // c9t259i25
	assign leaf[382] = !f[544] && !f[380] && f[488] && f[348]; // c9t259i25
	assign leaf[383] = !f[544] && f[380] && !f[467] && !f[412]; // c9t259i25
	assign leaf[384] = !f[544] && f[380] && !f[467] && f[412]; // c9t259i25
	assign leaf[385] = !f[544] && f[380] && f[467] && !f[356]; // c9t259i25
	assign leaf[386] = !f[544] && f[380] && f[467] && f[356]; // c9t259i25
	assign leaf[387] = f[544] && !f[629] && !f[488] && !f[273]; // c9t259i25
	assign leaf[388] = f[544] && !f[629] && !f[488] && f[273]; // c9t259i25
	assign leaf[389] = f[544] && !f[629] && f[488] && !f[399]; // c9t259i25
	assign leaf[390] = f[544] && !f[629] && f[488] && f[399]; // c9t259i25
	assign leaf[391] = f[544] && f[629] && !f[207] && !f[213]; // c9t259i25
	assign leaf[392] = f[544] && f[629] && !f[207] && f[213]; // c9t259i25
	assign leaf[393] = f[544] && f[629] && f[207] && !f[461]; // c9t259i25
	assign leaf[394] = f[544] && f[629] && f[207] && f[461]; // c9t259i25
	assign leaf[395] = !f[742] && !f[355] && !f[439] && !f[523]; // c9t269i26
	assign leaf[396] = !f[742] && !f[355] && !f[439] && f[523]; // c9t269i26
	assign leaf[397] = !f[742] && !f[355] && f[439] && !f[356]; // c9t269i26
	assign leaf[398] = !f[742] && !f[355] && f[439] && f[356]; // c9t269i26
	assign leaf[399] = !f[742] && f[355] && !f[213] && !f[318]; // c9t269i26
	assign leaf[400] = !f[742] && f[355] && !f[213] && f[318]; // c9t269i26
	assign leaf[401] = !f[742] && f[355] && f[213] && !f[566]; // c9t269i26
	assign leaf[402] = !f[742] && f[355] && f[213] && f[566]; // c9t269i26
	assign leaf[403] = f[742] && !f[323] && !f[488] && !f[406]; // c9t269i26
	assign leaf[404] = f[742] && !f[323] && !f[488] && f[406]; // c9t269i26
	assign leaf[405] = f[742] && !f[323] && f[488] && !f[546]; // c9t269i26
	assign leaf[406] = f[742] && !f[323] && f[488] && f[546]; // c9t269i26
	assign leaf[407] = f[742] && f[323] && !f[259] && !f[214]; // c9t269i26
	assign leaf[408] = f[742] && f[323] && !f[259] && f[214]; // c9t269i26
	assign leaf[409] = f[742] && f[323] && f[259] && !f[206]; // c9t269i26
	assign leaf[410] = f[742] && f[323] && f[259] && f[206]; // c9t269i26
	assign leaf[411] = !f[201] && !f[694] && !f[517] && !f[543]; // c9t279i27
	assign leaf[412] = !f[201] && !f[694] && !f[517] && f[543]; // c9t279i27
	assign leaf[413] = !f[201] && !f[694] && f[517] && !f[658]; // c9t279i27
	assign leaf[414] = !f[201] && !f[694] && f[517] && f[658]; // c9t279i27
	assign leaf[415] = !f[201] && f[694] && !f[403] && !f[666]; // c9t279i27
	assign leaf[416] = !f[201] && f[694] && !f[403] && f[666]; // c9t279i27
	assign leaf[417] = !f[201] && f[694] && f[403] && !f[313]; // c9t279i27
	assign leaf[418] = !f[201] && f[694] && f[403] && f[313]; // c9t279i27
	assign leaf[419] = f[201] && !f[379] && !f[665]; // c9t279i27
	assign leaf[420] = f[201] && !f[379] && f[665]; // c9t279i27
	assign leaf[421] = f[201] && f[379]; // c9t279i27
	assign leaf[422] = !f[594] && !f[129] && !f[149] && !f[379]; // c9t289i28
	assign leaf[423] = !f[594] && !f[129] && !f[149] && f[379]; // c9t289i28
	assign leaf[424] = !f[594] && !f[129] && f[149] && !f[258]; // c9t289i28
	assign leaf[425] = !f[594] && !f[129] && f[149] && f[258]; // c9t289i28
	assign leaf[426] = !f[594] && f[129] && !f[126]; // c9t289i28
	assign leaf[427] = !f[594] && f[129] && f[126] && !f[292]; // c9t289i28
	assign leaf[428] = !f[594] && f[129] && f[126] && f[292]; // c9t289i28
	assign leaf[429] = f[594] && !f[551] && !f[181]; // c9t289i28
	assign leaf[430] = f[594] && !f[551] && f[181] && !f[436]; // c9t289i28
	assign leaf[431] = f[594] && !f[551] && f[181] && f[436]; // c9t289i28
	assign leaf[432] = f[594] && f[551] && !f[399] && !f[211]; // c9t289i28
	assign leaf[433] = f[594] && f[551] && !f[399] && f[211]; // c9t289i28
	assign leaf[434] = f[594] && f[551] && f[399] && !f[466]; // c9t289i28
	assign leaf[435] = f[594] && f[551] && f[399] && f[466]; // c9t289i28
	assign leaf[436] = !f[342] && !f[495] && !f[319] && !f[317]; // c9t299i29
	assign leaf[437] = !f[342] && !f[495] && !f[319] && f[317]; // c9t299i29
	assign leaf[438] = !f[342] && !f[495] && f[319] && !f[379]; // c9t299i29
	assign leaf[439] = !f[342] && !f[495] && f[319] && f[379]; // c9t299i29
	assign leaf[440] = !f[342] && f[495] && !f[664] && !f[344]; // c9t299i29
	assign leaf[441] = !f[342] && f[495] && !f[664] && f[344]; // c9t299i29
	assign leaf[442] = !f[342] && f[495] && f[664] && !f[607]; // c9t299i29
	assign leaf[443] = !f[342] && f[495] && f[664] && f[607]; // c9t299i29
	assign leaf[444] = f[342] && !f[345] && !f[385] && !f[213]; // c9t299i29
	assign leaf[445] = f[342] && !f[345] && !f[385] && f[213]; // c9t299i29
	assign leaf[446] = f[342] && !f[345] && f[385] && !f[343]; // c9t299i29
	assign leaf[447] = f[342] && !f[345] && f[385] && f[343]; // c9t299i29
	assign leaf[448] = f[342] && f[345] && !f[456] && !f[206]; // c9t299i29
	assign leaf[449] = f[342] && f[345] && !f[456] && f[206]; // c9t299i29
	assign leaf[450] = f[342] && f[345] && f[456] && !f[410]; // c9t299i29
	assign leaf[451] = f[342] && f[345] && f[456] && f[410]; // c9t299i29
	assign leaf[452] = !f[161] && !f[572] && !f[188] && !f[209]; // c9t309i30
	assign leaf[453] = !f[161] && !f[572] && !f[188] && f[209]; // c9t309i30
	assign leaf[454] = !f[161] && !f[572] && f[188] && !f[601]; // c9t309i30
	assign leaf[455] = !f[161] && !f[572] && f[188] && f[601]; // c9t309i30
	assign leaf[456] = !f[161] && f[572] && !f[207] && !f[214]; // c9t309i30
	assign leaf[457] = !f[161] && f[572] && !f[207] && f[214]; // c9t309i30
	assign leaf[458] = !f[161] && f[572] && f[207] && !f[461]; // c9t309i30
	assign leaf[459] = !f[161] && f[572] && f[207] && f[461]; // c9t309i30
	assign leaf[460] = f[161] && !f[329]; // c9t309i30
	assign leaf[461] = f[161] && f[329] && !f[601] && !f[319]; // c9t309i30
	assign leaf[462] = f[161] && f[329] && !f[601] && f[319]; // c9t309i30
	assign leaf[463] = f[161] && f[329] && f[601]; // c9t309i30
	assign leaf[464] = !f[631] && !f[715] && !f[566] && !f[350]; // c9t319i31
	assign leaf[465] = !f[631] && !f[715] && !f[566] && f[350]; // c9t319i31
	assign leaf[466] = !f[631] && !f[715] && f[566] && !f[606]; // c9t319i31
	assign leaf[467] = !f[631] && !f[715] && f[566] && f[606]; // c9t319i31
	assign leaf[468] = !f[631] && f[715] && !f[381] && !f[294]; // c9t319i31
	assign leaf[469] = !f[631] && f[715] && !f[381] && f[294]; // c9t319i31
	assign leaf[470] = !f[631] && f[715] && f[381] && !f[743]; // c9t319i31
	assign leaf[471] = !f[631] && f[715] && f[381] && f[743]; // c9t319i31
	assign leaf[472] = f[631] && !f[545] && !f[209] && !f[742]; // c9t319i31
	assign leaf[473] = f[631] && !f[545] && !f[209] && f[742]; // c9t319i31
	assign leaf[474] = f[631] && !f[545] && f[209] && !f[237]; // c9t319i31
	assign leaf[475] = f[631] && !f[545] && f[209] && f[237]; // c9t319i31
	assign leaf[476] = f[631] && f[545] && !f[485] && !f[489]; // c9t319i31
	assign leaf[477] = f[631] && f[545] && !f[485] && f[489]; // c9t319i31
	assign leaf[478] = f[631] && f[545] && f[485] && !f[576]; // c9t319i31
	assign leaf[479] = f[631] && f[545] && f[485] && f[576]; // c9t319i31
	assign leaf[480] = !f[693] && !f[608] && !f[351] && !f[385]; // c9t329i32
	assign leaf[481] = !f[693] && !f[608] && !f[351] && f[385]; // c9t329i32
	assign leaf[482] = !f[693] && !f[608] && f[351] && !f[461]; // c9t329i32
	assign leaf[483] = !f[693] && !f[608] && f[351] && f[461]; // c9t329i32
	assign leaf[484] = !f[693] && f[608] && !f[692] && !f[330]; // c9t329i32
	assign leaf[485] = !f[693] && f[608] && !f[692] && f[330]; // c9t329i32
	assign leaf[486] = !f[693] && f[608] && f[692] && !f[318]; // c9t329i32
	assign leaf[487] = !f[693] && f[608] && f[692] && f[318]; // c9t329i32
	assign leaf[488] = f[693] && !f[229] && !f[320] && !f[203]; // c9t329i32
	assign leaf[489] = f[693] && !f[229] && !f[320] && f[203]; // c9t329i32
	assign leaf[490] = f[693] && !f[229] && f[320] && !f[461]; // c9t329i32
	assign leaf[491] = f[693] && !f[229] && f[320] && f[461]; // c9t329i32
	assign leaf[492] = f[693] && f[229] && !f[429]; // c9t329i32
	assign leaf[493] = f[693] && f[229] && f[429] && !f[407]; // c9t329i32
	assign leaf[494] = f[693] && f[229] && f[429] && f[407]; // c9t329i32
	assign leaf[495] = !f[436] && !f[465] && !f[667] && !f[492]; // c9t339i33
	assign leaf[496] = !f[436] && !f[465] && !f[667] && f[492]; // c9t339i33
	assign leaf[497] = !f[436] && !f[465] && f[667] && !f[454]; // c9t339i33
	assign leaf[498] = !f[436] && !f[465] && f[667] && f[454]; // c9t339i33
	assign leaf[499] = !f[436] && f[465] && !f[293] && !f[462]; // c9t339i33
	assign leaf[500] = !f[436] && f[465] && !f[293] && f[462]; // c9t339i33
	assign leaf[501] = !f[436] && f[465] && f[293] && !f[433]; // c9t339i33
	assign leaf[502] = !f[436] && f[465] && f[293] && f[433]; // c9t339i33
	assign leaf[503] = f[436] && !f[469] && !f[572] && !f[413]; // c9t339i33
	assign leaf[504] = f[436] && !f[469] && !f[572] && f[413]; // c9t339i33
	assign leaf[505] = f[436] && !f[469] && f[572] && !f[346]; // c9t339i33
	assign leaf[506] = f[436] && !f[469] && f[572] && f[346]; // c9t339i33
	assign leaf[507] = f[436] && f[469] && !f[357] && !f[692]; // c9t339i33
	assign leaf[508] = f[436] && f[469] && !f[357] && f[692]; // c9t339i33
	assign leaf[509] = f[436] && f[469] && f[357] && !f[347]; // c9t339i33
	assign leaf[510] = f[436] && f[469] && f[357] && f[347]; // c9t339i33
	assign leaf[511] = !f[229] && !f[162] && !f[175] && !f[639]; // c9t349i34
	assign leaf[512] = !f[229] && !f[162] && !f[175] && f[639]; // c9t349i34
	assign leaf[513] = !f[229] && !f[162] && f[175] && !f[151]; // c9t349i34
	assign leaf[514] = !f[229] && !f[162] && f[175] && f[151]; // c9t349i34
	assign leaf[515] = !f[229] && f[162] && !f[679]; // c9t349i34
	assign leaf[516] = !f[229] && f[162] && f[679]; // c9t349i34
	assign leaf[517] = f[229] && !f[151] && !f[407] && !f[429]; // c9t349i34
	assign leaf[518] = f[229] && !f[151] && !f[407] && f[429]; // c9t349i34
	assign leaf[519] = f[229] && !f[151] && f[407]; // c9t349i34
	assign leaf[520] = f[229] && f[151]; // c9t349i34
	assign leaf[521] = !f[742] && !f[632] && !f[688] && !f[542]; // c9t359i35
	assign leaf[522] = !f[742] && !f[632] && !f[688] && f[542]; // c9t359i35
	assign leaf[523] = !f[742] && !f[632] && f[688] && !f[662]; // c9t359i35
	assign leaf[524] = !f[742] && !f[632] && f[688] && f[662]; // c9t359i35
	assign leaf[525] = !f[742] && f[632] && !f[493] && !f[517]; // c9t359i35
	assign leaf[526] = !f[742] && f[632] && !f[493] && f[517]; // c9t359i35
	assign leaf[527] = !f[742] && f[632] && f[493] && !f[182]; // c9t359i35
	assign leaf[528] = !f[742] && f[632] && f[493] && f[182]; // c9t359i35
	assign leaf[529] = f[742] && !f[634] && !f[204] && !f[290]; // c9t359i35
	assign leaf[530] = f[742] && !f[634] && !f[204] && f[290]; // c9t359i35
	assign leaf[531] = f[742] && !f[634] && f[204]; // c9t359i35
	assign leaf[532] = f[742] && f[634]; // c9t359i35
	assign leaf[533] = !f[356] && !f[468] && !f[412] && !f[244]; // c9t369i36
	assign leaf[534] = !f[356] && !f[468] && !f[412] && f[244]; // c9t369i36
	assign leaf[535] = !f[356] && !f[468] && f[412] && !f[495]; // c9t369i36
	assign leaf[536] = !f[356] && !f[468] && f[412] && f[495]; // c9t369i36
	assign leaf[537] = !f[356] && f[468] && !f[408] && !f[287]; // c9t369i36
	assign leaf[538] = !f[356] && f[468] && !f[408] && f[287]; // c9t369i36
	assign leaf[539] = !f[356] && f[468] && f[408] && !f[694]; // c9t369i36
	assign leaf[540] = !f[356] && f[468] && f[408] && f[694]; // c9t369i36
	assign leaf[541] = f[356] && !f[411] && !f[741] && !f[437]; // c9t369i36
	assign leaf[542] = f[356] && !f[411] && !f[741] && f[437]; // c9t369i36
	assign leaf[543] = f[356] && !f[411] && f[741]; // c9t369i36
	assign leaf[544] = f[356] && f[411] && !f[213] && !f[185]; // c9t369i36
	assign leaf[545] = f[356] && f[411] && !f[213] && f[185]; // c9t369i36
	assign leaf[546] = f[356] && f[411] && f[213] && !f[295]; // c9t369i36
	assign leaf[547] = f[356] && f[411] && f[213] && f[295]; // c9t369i36
	assign leaf[548] = !f[191] && !f[319] && !f[371] && !f[345]; // c9t379i37
	assign leaf[549] = !f[191] && !f[319] && !f[371] && f[345]; // c9t379i37
	assign leaf[550] = !f[191] && !f[319] && f[371] && !f[345]; // c9t379i37
	assign leaf[551] = !f[191] && !f[319] && f[371] && f[345]; // c9t379i37
	assign leaf[552] = !f[191] && f[319] && !f[522] && !f[467]; // c9t379i37
	assign leaf[553] = !f[191] && f[319] && !f[522] && f[467]; // c9t379i37
	assign leaf[554] = !f[191] && f[319] && f[522] && !f[410]; // c9t379i37
	assign leaf[555] = !f[191] && f[319] && f[522] && f[410]; // c9t379i37
	assign leaf[556] = f[191] && !f[273] && !f[399]; // c9t379i37
	assign leaf[557] = f[191] && !f[273] && f[399]; // c9t379i37
	assign leaf[558] = f[191] && f[273] && !f[482]; // c9t379i37
	assign leaf[559] = f[191] && f[273] && f[482]; // c9t379i37
	assign leaf[560] = !f[368] && !f[437] && !f[549] && !f[382]; // c9t389i38
	assign leaf[561] = !f[368] && !f[437] && !f[549] && f[382]; // c9t389i38
	assign leaf[562] = !f[368] && !f[437] && f[549] && !f[462]; // c9t389i38
	assign leaf[563] = !f[368] && !f[437] && f[549] && f[462]; // c9t389i38
	assign leaf[564] = !f[368] && f[437] && !f[496] && !f[441]; // c9t389i38
	assign leaf[565] = !f[368] && f[437] && !f[496] && f[441]; // c9t389i38
	assign leaf[566] = !f[368] && f[437] && f[496] && !f[412]; // c9t389i38
	assign leaf[567] = !f[368] && f[437] && f[496] && f[412]; // c9t389i38
	assign leaf[568] = f[368] && !f[373] && !f[349] && !f[354]; // c9t389i38
	assign leaf[569] = f[368] && !f[373] && !f[349] && f[354]; // c9t389i38
	assign leaf[570] = f[368] && !f[373] && f[349]; // c9t389i38
	assign leaf[571] = f[368] && f[373] && !f[465]; // c9t389i38
	assign leaf[572] = f[368] && f[373] && f[465] && !f[260]; // c9t389i38
	assign leaf[573] = f[368] && f[373] && f[465] && f[260]; // c9t389i38
	assign leaf[574] = !f[350] && !f[486] && !f[406] && !f[512]; // c9t399i39
	assign leaf[575] = !f[350] && !f[486] && !f[406] && f[512]; // c9t399i39
	assign leaf[576] = !f[350] && !f[486] && f[406] && !f[489]; // c9t399i39
	assign leaf[577] = !f[350] && !f[486] && f[406] && f[489]; // c9t399i39
	assign leaf[578] = !f[350] && f[486] && !f[431] && !f[428]; // c9t399i39
	assign leaf[579] = !f[350] && f[486] && !f[431] && f[428]; // c9t399i39
	assign leaf[580] = !f[350] && f[486] && f[431] && !f[428]; // c9t399i39
	assign leaf[581] = !f[350] && f[486] && f[431] && f[428]; // c9t399i39
	assign leaf[582] = f[350] && !f[325] && !f[434] && !f[464]; // c9t399i39
	assign leaf[583] = f[350] && !f[325] && !f[434] && f[464]; // c9t399i39
	assign leaf[584] = f[350] && !f[325] && f[434] && !f[264]; // c9t399i39
	assign leaf[585] = f[350] && !f[325] && f[434] && f[264]; // c9t399i39
	assign leaf[586] = f[350] && f[325] && !f[460] && !f[456]; // c9t399i39
	assign leaf[587] = f[350] && f[325] && !f[460] && f[456]; // c9t399i39
	assign leaf[588] = f[350] && f[325] && f[460] && !f[345]; // c9t399i39
	assign leaf[589] = f[350] && f[325] && f[460] && f[345]; // c9t399i39
	assign leaf[590] = !f[408] && !f[439] && !f[410] && !f[550]; // c9t409i40
	assign leaf[591] = !f[408] && !f[439] && !f[410] && f[550]; // c9t409i40
	assign leaf[592] = !f[408] && !f[439] && f[410] && !f[324]; // c9t409i40
	assign leaf[593] = !f[408] && !f[439] && f[410] && f[324]; // c9t409i40
	assign leaf[594] = !f[408] && f[439] && !f[373] && !f[207]; // c9t409i40
	assign leaf[595] = !f[408] && f[439] && !f[373] && f[207]; // c9t409i40
	assign leaf[596] = !f[408] && f[439] && f[373] && !f[155]; // c9t409i40
	assign leaf[597] = !f[408] && f[439] && f[373] && f[155]; // c9t409i40
	assign leaf[598] = f[408] && !f[149] && !f[517] && !f[181]; // c9t409i40
	assign leaf[599] = f[408] && !f[149] && !f[517] && f[181]; // c9t409i40
	assign leaf[600] = f[408] && !f[149] && f[517] && !f[630]; // c9t409i40
	assign leaf[601] = f[408] && !f[149] && f[517] && f[630]; // c9t409i40
	assign leaf[602] = f[408] && f[149] && !f[286]; // c9t409i40
	assign leaf[603] = f[408] && f[149] && f[286]; // c9t409i40
	assign leaf[604] = !f[500] && !f[273] && !f[327] && !f[439]; // c9t419i41
	assign leaf[605] = !f[500] && !f[273] && !f[327] && f[439]; // c9t419i41
	assign leaf[606] = !f[500] && !f[273] && f[327] && !f[351]; // c9t419i41
	assign leaf[607] = !f[500] && !f[273] && f[327] && f[351]; // c9t419i41
	assign leaf[608] = !f[500] && f[273] && !f[215] && !f[241]; // c9t419i41
	assign leaf[609] = !f[500] && f[273] && !f[215] && f[241]; // c9t419i41
	assign leaf[610] = !f[500] && f[273] && f[215] && !f[385]; // c9t419i41
	assign leaf[611] = !f[500] && f[273] && f[215] && f[385]; // c9t419i41
	assign leaf[612] = f[500] && !f[416]; // c9t419i41
	assign leaf[613] = f[500] && f[416]; // c9t419i41
	assign leaf[614] = !f[350] && !f[406] && !f[487] && !f[514]; // c9t429i42
	assign leaf[615] = !f[350] && !f[406] && !f[487] && f[514]; // c9t429i42
	assign leaf[616] = !f[350] && !f[406] && f[487] && !f[404]; // c9t429i42
	assign leaf[617] = !f[350] && !f[406] && f[487] && f[404]; // c9t429i42
	assign leaf[618] = !f[350] && f[406] && !f[292] && !f[462]; // c9t429i42
	assign leaf[619] = !f[350] && f[406] && !f[292] && f[462]; // c9t429i42
	assign leaf[620] = !f[350] && f[406] && f[292] && !f[181]; // c9t429i42
	assign leaf[621] = !f[350] && f[406] && f[292] && f[181]; // c9t429i42
	assign leaf[622] = f[350] && !f[487] && !f[324] && !f[608]; // c9t429i42
	assign leaf[623] = f[350] && !f[487] && !f[324] && f[608]; // c9t429i42
	assign leaf[624] = f[350] && !f[487] && f[324] && !f[461]; // c9t429i42
	assign leaf[625] = f[350] && !f[487] && f[324] && f[461]; // c9t429i42
	assign leaf[626] = f[350] && f[487] && !f[434] && !f[580]; // c9t429i42
	assign leaf[627] = f[350] && f[487] && !f[434] && f[580]; // c9t429i42
	assign leaf[628] = f[350] && f[487] && f[434] && !f[600]; // c9t429i42
	assign leaf[629] = f[350] && f[487] && f[434] && f[600]; // c9t429i42
	assign leaf[630] = !f[472] && !f[201] && !f[315] && !f[205]; // c9t439i43
	assign leaf[631] = !f[472] && !f[201] && !f[315] && f[205]; // c9t439i43
	assign leaf[632] = !f[472] && !f[201] && f[315] && !f[317]; // c9t439i43
	assign leaf[633] = !f[472] && !f[201] && f[315] && f[317]; // c9t439i43
	assign leaf[634] = !f[472] && f[201] && !f[666]; // c9t439i43
	assign leaf[635] = !f[472] && f[201] && f[666]; // c9t439i43
	assign leaf[636] = f[472]; // c9t439i43
	assign leaf[637] = !f[740] && !f[742] && !f[709] && !f[182]; // c9t449i44
	assign leaf[638] = !f[740] && !f[742] && !f[709] && f[182]; // c9t449i44
	assign leaf[639] = !f[740] && !f[742] && f[709] && !f[236]; // c9t449i44
	assign leaf[640] = !f[740] && !f[742] && f[709] && f[236]; // c9t449i44
	assign leaf[641] = !f[740] && f[742] && !f[242] && !f[268]; // c9t449i44
	assign leaf[642] = !f[740] && f[742] && !f[242] && f[268]; // c9t449i44
	assign leaf[643] = !f[740] && f[742] && f[242] && !f[206]; // c9t449i44
	assign leaf[644] = !f[740] && f[742] && f[242] && f[206]; // c9t449i44
	assign leaf[645] = f[740] && !f[243] && !f[406] && !f[711]; // c9t449i44
	assign leaf[646] = f[740] && !f[243] && !f[406] && f[711]; // c9t449i44
	assign leaf[647] = f[740] && !f[243] && f[406] && !f[377]; // c9t449i44
	assign leaf[648] = f[740] && !f[243] && f[406] && f[377]; // c9t449i44
	assign leaf[649] = f[740] && f[243] && !f[235] && !f[404]; // c9t449i44
	assign leaf[650] = f[740] && f[243] && !f[235] && f[404]; // c9t449i44
	assign leaf[651] = f[740] && f[243] && f[235] && !f[349]; // c9t449i44
	assign leaf[652] = f[740] && f[243] && f[235] && f[349]; // c9t449i44
	assign leaf[653] = !f[746] && !f[734] && !f[275] && !f[606]; // c9t459i45
	assign leaf[654] = !f[746] && !f[734] && !f[275] && f[606]; // c9t459i45
	assign leaf[655] = !f[746] && !f[734] && f[275] && !f[215]; // c9t459i45
	assign leaf[656] = !f[746] && !f[734] && f[275] && f[215]; // c9t459i45
	assign leaf[657] = !f[746] && f[734] && !f[431]; // c9t459i45
	assign leaf[658] = !f[746] && f[734] && f[431]; // c9t459i45
	assign leaf[659] = f[746] && !f[431] && !f[291] && !f[243]; // c9t459i45
	assign leaf[660] = f[746] && !f[431] && !f[291] && f[243]; // c9t459i45
	assign leaf[661] = f[746] && !f[431] && f[291] && !f[401]; // c9t459i45
	assign leaf[662] = f[746] && !f[431] && f[291] && f[401]; // c9t459i45
	assign leaf[663] = f[746] && f[431] && !f[661]; // c9t459i45
	assign leaf[664] = f[746] && f[431] && f[661]; // c9t459i45
	assign leaf[665] = !f[368] && !f[415] && !f[353] && !f[405]; // c9t469i46
	assign leaf[666] = !f[368] && !f[415] && !f[353] && f[405]; // c9t469i46
	assign leaf[667] = !f[368] && !f[415] && f[353] && !f[378]; // c9t469i46
	assign leaf[668] = !f[368] && !f[415] && f[353] && f[378]; // c9t469i46
	assign leaf[669] = !f[368] && f[415] && !f[313] && !f[682]; // c9t469i46
	assign leaf[670] = !f[368] && f[415] && !f[313] && f[682]; // c9t469i46
	assign leaf[671] = !f[368] && f[415] && f[313]; // c9t469i46
	assign leaf[672] = f[368] && !f[373] && !f[660] && !f[326]; // c9t469i46
	assign leaf[673] = f[368] && !f[373] && !f[660] && f[326]; // c9t469i46
	assign leaf[674] = f[368] && !f[373] && f[660] && !f[434]; // c9t469i46
	assign leaf[675] = f[368] && !f[373] && f[660] && f[434]; // c9t469i46
	assign leaf[676] = f[368] && f[373] && !f[286]; // c9t469i46
	assign leaf[677] = f[368] && f[373] && f[286] && !f[238]; // c9t469i46
	assign leaf[678] = f[368] && f[373] && f[286] && f[238]; // c9t469i46
	assign leaf[679] = !f[274] && !f[356] && !f[323] && !f[523]; // c9t479i47
	assign leaf[680] = !f[274] && !f[356] && !f[323] && f[523]; // c9t479i47
	assign leaf[681] = !f[274] && !f[356] && f[323] && !f[434]; // c9t479i47
	assign leaf[682] = !f[274] && !f[356] && f[323] && f[434]; // c9t479i47
	assign leaf[683] = !f[274] && f[356] && !f[466] && !f[328]; // c9t479i47
	assign leaf[684] = !f[274] && f[356] && !f[466] && f[328]; // c9t479i47
	assign leaf[685] = !f[274] && f[356] && f[466] && !f[128]; // c9t479i47
	assign leaf[686] = !f[274] && f[356] && f[466] && f[128]; // c9t479i47
	assign leaf[687] = f[274] && !f[215] && !f[242] && !f[158]; // c9t479i47
	assign leaf[688] = f[274] && !f[215] && !f[242] && f[158]; // c9t479i47
	assign leaf[689] = f[274] && !f[215] && f[242] && !f[375]; // c9t479i47
	assign leaf[690] = f[274] && !f[215] && f[242] && f[375]; // c9t479i47
	assign leaf[691] = f[274] && f[215] && !f[211] && !f[408]; // c9t479i47
	assign leaf[692] = f[274] && f[215] && !f[211] && f[408]; // c9t479i47
	assign leaf[693] = f[274] && f[215] && f[211] && !f[412]; // c9t479i47
	assign leaf[694] = f[274] && f[215] && f[211] && f[412]; // c9t479i47
	assign leaf[695] = !f[162] && !f[175] && !f[229] && !f[720]; // c9t489i48
	assign leaf[696] = !f[162] && !f[175] && !f[229] && f[720]; // c9t489i48
	assign leaf[697] = !f[162] && !f[175] && f[229] && !f[369]; // c9t489i48
	assign leaf[698] = !f[162] && !f[175] && f[229] && f[369]; // c9t489i48
	assign leaf[699] = !f[162] && f[175] && !f[257] && !f[353]; // c9t489i48
	assign leaf[700] = !f[162] && f[175] && !f[257] && f[353]; // c9t489i48
	assign leaf[701] = !f[162] && f[175] && f[257] && !f[266]; // c9t489i48
	assign leaf[702] = !f[162] && f[175] && f[257] && f[266]; // c9t489i48
	assign leaf[703] = f[162]; // c9t489i48
	assign leaf[704] = !f[573] && !f[711] && !f[404] && !f[461]; // c9t499i49
	assign leaf[705] = !f[573] && !f[711] && !f[404] && f[461]; // c9t499i49
	assign leaf[706] = !f[573] && !f[711] && f[404] && !f[456]; // c9t499i49
	assign leaf[707] = !f[573] && !f[711] && f[404] && f[456]; // c9t499i49
	assign leaf[708] = !f[573] && f[711] && !f[412] && !f[600]; // c9t499i49
	assign leaf[709] = !f[573] && f[711] && !f[412] && f[600]; // c9t499i49
	assign leaf[710] = !f[573] && f[711] && f[412] && !f[494]; // c9t499i49
	assign leaf[711] = !f[573] && f[711] && f[412] && f[494]; // c9t499i49
	assign leaf[712] = f[573] && !f[207] && !f[549] && !f[489]; // c9t499i49
	assign leaf[713] = f[573] && !f[207] && !f[549] && f[489]; // c9t499i49
	assign leaf[714] = f[573] && !f[207] && f[549] && !f[484]; // c9t499i49
	assign leaf[715] = f[573] && !f[207] && f[549] && f[484]; // c9t499i49
	assign leaf[716] = f[573] && f[207] && !f[489] && !f[458]; // c9t499i49
	assign leaf[717] = f[573] && f[207] && !f[489] && f[458]; // c9t499i49
	assign leaf[718] = f[573] && f[207] && f[489] && !f[290]; // c9t499i49
	assign leaf[719] = f[573] && f[207] && f[489] && f[290]; // c9t499i49
	assign leaf[720] = !f[129] && !f[415] && !f[244] && !f[326]; // c9t509i50
	assign leaf[721] = !f[129] && !f[415] && !f[244] && f[326]; // c9t509i50
	assign leaf[722] = !f[129] && !f[415] && f[244] && !f[330]; // c9t509i50
	assign leaf[723] = !f[129] && !f[415] && f[244] && f[330]; // c9t509i50
	assign leaf[724] = !f[129] && f[415] && !f[302] && !f[430]; // c9t509i50
	assign leaf[725] = !f[129] && f[415] && !f[302] && f[430]; // c9t509i50
	assign leaf[726] = !f[129] && f[415] && f[302] && !f[403]; // c9t509i50
	assign leaf[727] = !f[129] && f[415] && f[302] && f[403]; // c9t509i50
	assign leaf[728] = f[129] && !f[217] && !f[185]; // c9t509i50
	assign leaf[729] = f[129] && !f[217] && f[185]; // c9t509i50
	assign leaf[730] = f[129] && f[217]; // c9t509i50
	assign leaf[731] = !f[340] && !f[353] && !f[385] && !f[156]; // c9t519i51
	assign leaf[732] = !f[340] && !f[353] && !f[385] && f[156]; // c9t519i51
	assign leaf[733] = !f[340] && !f[353] && f[385] && !f[214]; // c9t519i51
	assign leaf[734] = !f[340] && !f[353] && f[385] && f[214]; // c9t519i51
	assign leaf[735] = !f[340] && f[353] && !f[574] && !f[712]; // c9t519i51
	assign leaf[736] = !f[340] && f[353] && !f[574] && f[712]; // c9t519i51
	assign leaf[737] = !f[340] && f[353] && f[574] && !f[543]; // c9t519i51
	assign leaf[738] = !f[340] && f[353] && f[574] && f[543]; // c9t519i51
	assign leaf[739] = f[340] && !f[346] && !f[688] && !f[526]; // c9t519i51
	assign leaf[740] = f[340] && !f[346] && !f[688] && f[526]; // c9t519i51
	assign leaf[741] = f[340] && !f[346] && f[688]; // c9t519i51
	assign leaf[742] = f[340] && f[346] && !f[214]; // c9t519i51
	assign leaf[743] = f[340] && f[346] && f[214]; // c9t519i51
	assign leaf[744] = !f[584] && !f[500] && !f[740] && !f[326]; // c9t529i52
	assign leaf[745] = !f[584] && !f[500] && !f[740] && f[326]; // c9t529i52
	assign leaf[746] = !f[584] && !f[500] && f[740] && !f[714]; // c9t529i52
	assign leaf[747] = !f[584] && !f[500] && f[740] && f[714]; // c9t529i52
	assign leaf[748] = !f[584] && f[500]; // c9t529i52
	assign leaf[749] = f[584] && !f[297]; // c9t529i52
	assign leaf[750] = f[584] && f[297]; // c9t529i52
	assign leaf[751] = !f[605] && !f[566] && !f[717] && !f[378]; // c9t539i53
	assign leaf[752] = !f[605] && !f[566] && !f[717] && f[378]; // c9t539i53
	assign leaf[753] = !f[605] && !f[566] && f[717] && !f[233]; // c9t539i53
	assign leaf[754] = !f[605] && !f[566] && f[717] && f[233]; // c9t539i53
	assign leaf[755] = !f[605] && f[566] && !f[631]; // c9t539i53
	assign leaf[756] = !f[605] && f[566] && f[631]; // c9t539i53
	assign leaf[757] = f[605] && !f[546] && !f[180] && !f[236]; // c9t539i53
	assign leaf[758] = f[605] && !f[546] && !f[180] && f[236]; // c9t539i53
	assign leaf[759] = f[605] && !f[546] && f[180] && !f[265]; // c9t539i53
	assign leaf[760] = f[605] && !f[546] && f[180] && f[265]; // c9t539i53
	assign leaf[761] = f[605] && f[546] && !f[494] && !f[512]; // c9t539i53
	assign leaf[762] = f[605] && f[546] && !f[494] && f[512]; // c9t539i53
	assign leaf[763] = f[605] && f[546] && f[494] && !f[469]; // c9t539i53
	assign leaf[764] = f[605] && f[546] && f[494] && f[469]; // c9t539i53
	assign leaf[765] = !f[323] && !f[355] && !f[297] && !f[463]; // c9t549i54
	assign leaf[766] = !f[323] && !f[355] && !f[297] && f[463]; // c9t549i54
	assign leaf[767] = !f[323] && !f[355] && f[297] && !f[241]; // c9t549i54
	assign leaf[768] = !f[323] && !f[355] && f[297] && f[241]; // c9t549i54
	assign leaf[769] = !f[323] && f[355] && !f[407] && !f[515]; // c9t549i54
	assign leaf[770] = !f[323] && f[355] && !f[407] && f[515]; // c9t549i54
	assign leaf[771] = !f[323] && f[355] && f[407] && !f[213]; // c9t549i54
	assign leaf[772] = !f[323] && f[355] && f[407] && f[213]; // c9t549i54
	assign leaf[773] = f[323] && !f[295] && !f[188] && !f[519]; // c9t549i54
	assign leaf[774] = f[323] && !f[295] && !f[188] && f[519]; // c9t549i54
	assign leaf[775] = f[323] && !f[295] && f[188] && !f[683]; // c9t549i54
	assign leaf[776] = f[323] && !f[295] && f[188] && f[683]; // c9t549i54
	assign leaf[777] = f[323] && f[295] && !f[575] && !f[179]; // c9t549i54
	assign leaf[778] = f[323] && f[295] && !f[575] && f[179]; // c9t549i54
	assign leaf[779] = f[323] && f[295] && f[575] && !f[489]; // c9t549i54
	assign leaf[780] = f[323] && f[295] && f[575] && f[489]; // c9t549i54
	assign leaf[781] = !f[742] && !f[686] && !f[740] && !f[602]; // c9t559i55
	assign leaf[782] = !f[742] && !f[686] && !f[740] && f[602]; // c9t559i55
	assign leaf[783] = !f[742] && !f[686] && f[740] && !f[710]; // c9t559i55
	assign leaf[784] = !f[742] && !f[686] && f[740] && f[710]; // c9t559i55
	assign leaf[785] = !f[742] && f[686] && !f[545] && !f[408]; // c9t559i55
	assign leaf[786] = !f[742] && f[686] && !f[545] && f[408]; // c9t559i55
	assign leaf[787] = !f[742] && f[686] && f[545] && !f[184]; // c9t559i55
	assign leaf[788] = !f[742] && f[686] && f[545] && f[184]; // c9t559i55
	assign leaf[789] = f[742] && !f[242] && !f[405] && !f[322]; // c9t559i55
	assign leaf[790] = f[742] && !f[242] && !f[405] && f[322]; // c9t559i55
	assign leaf[791] = f[742] && !f[242] && f[405] && !f[326]; // c9t559i55
	assign leaf[792] = f[742] && !f[242] && f[405] && f[326]; // c9t559i55
	assign leaf[793] = f[742] && f[242] && !f[684] && !f[488]; // c9t559i55
	assign leaf[794] = f[742] && f[242] && !f[684] && f[488]; // c9t559i55
	assign leaf[795] = f[742] && f[242] && f[684]; // c9t559i55
	assign leaf[796] = !f[131] && !f[369] && !f[441] && !f[497]; // c9t569i56
	assign leaf[797] = !f[131] && !f[369] && !f[441] && f[497]; // c9t569i56
	assign leaf[798] = !f[131] && !f[369] && f[441] && !f[544]; // c9t569i56
	assign leaf[799] = !f[131] && !f[369] && f[441] && f[544]; // c9t569i56
	assign leaf[800] = !f[131] && f[369] && !f[346] && !f[359]; // c9t569i56
	assign leaf[801] = !f[131] && f[369] && !f[346] && f[359]; // c9t569i56
	assign leaf[802] = !f[131] && f[369] && f[346] && !f[386]; // c9t569i56
	assign leaf[803] = !f[131] && f[369] && f[346] && f[386]; // c9t569i56
	assign leaf[804] = f[131] && !f[509]; // c9t569i56
	assign leaf[805] = f[131] && f[509]; // c9t569i56
	assign leaf[806] = !f[734] && !f[380] && !f[440] && !f[325]; // c9t579i57
	assign leaf[807] = !f[734] && !f[380] && !f[440] && f[325]; // c9t579i57
	assign leaf[808] = !f[734] && !f[380] && f[440] && !f[543]; // c9t579i57
	assign leaf[809] = !f[734] && !f[380] && f[440] && f[543]; // c9t579i57
	assign leaf[810] = !f[734] && f[380] && !f[467] && !f[523]; // c9t579i57
	assign leaf[811] = !f[734] && f[380] && !f[467] && f[523]; // c9t579i57
	assign leaf[812] = !f[734] && f[380] && f[467] && !f[343]; // c9t579i57
	assign leaf[813] = !f[734] && f[380] && f[467] && f[343]; // c9t579i57
	assign leaf[814] = f[734] && !f[597]; // c9t579i57
	assign leaf[815] = f[734] && f[597]; // c9t579i57
	assign leaf[816] = !f[149] && !f[388] && !f[508] && !f[256]; // c9t589i58
	assign leaf[817] = !f[149] && !f[388] && !f[508] && f[256]; // c9t589i58
	assign leaf[818] = !f[149] && !f[388] && f[508] && !f[662]; // c9t589i58
	assign leaf[819] = !f[149] && !f[388] && f[508] && f[662]; // c9t589i58
	assign leaf[820] = !f[149] && f[388]; // c9t589i58
	assign leaf[821] = f[149] && !f[286]; // c9t589i58
	assign leaf[822] = f[149] && f[286] && !f[354]; // c9t589i58
	assign leaf[823] = f[149] && f[286] && f[354]; // c9t589i58
	assign leaf[824] = !f[131] && !f[178] && !f[259] && !f[205]; // c9t599i59
	assign leaf[825] = !f[131] && !f[178] && !f[259] && f[205]; // c9t599i59
	assign leaf[826] = !f[131] && !f[178] && f[259] && !f[206]; // c9t599i59
	assign leaf[827] = !f[131] && !f[178] && f[259] && f[206]; // c9t599i59
	assign leaf[828] = !f[131] && f[178] && !f[181] && !f[691]; // c9t599i59
	assign leaf[829] = !f[131] && f[178] && !f[181] && f[691]; // c9t599i59
	assign leaf[830] = !f[131] && f[178] && f[181] && !f[210]; // c9t599i59
	assign leaf[831] = !f[131] && f[178] && f[181] && f[210]; // c9t599i59
	assign leaf[832] = f[131] && !f[128]; // c9t599i59
	assign leaf[833] = f[131] && f[128]; // c9t599i59
	assign leaf[834] = !f[709] && !f[627] && !f[404] && !f[182]; // c9t609i60
	assign leaf[835] = !f[709] && !f[627] && !f[404] && f[182]; // c9t609i60
	assign leaf[836] = !f[709] && !f[627] && f[404] && !f[378]; // c9t609i60
	assign leaf[837] = !f[709] && !f[627] && f[404] && f[378]; // c9t609i60
	assign leaf[838] = !f[709] && f[627] && !f[516] && !f[485]; // c9t609i60
	assign leaf[839] = !f[709] && f[627] && !f[516] && f[485]; // c9t609i60
	assign leaf[840] = !f[709] && f[627] && f[516] && !f[186]; // c9t609i60
	assign leaf[841] = !f[709] && f[627] && f[516] && f[186]; // c9t609i60
	assign leaf[842] = f[709] && !f[264] && !f[293] && !f[316]; // c9t609i60
	assign leaf[843] = f[709] && !f[264] && !f[293] && f[316]; // c9t609i60
	assign leaf[844] = f[709] && !f[264] && f[293] && !f[375]; // c9t609i60
	assign leaf[845] = f[709] && !f[264] && f[293] && f[375]; // c9t609i60
	assign leaf[846] = f[709] && f[264] && !f[213] && !f[268]; // c9t609i60
	assign leaf[847] = f[709] && f[264] && !f[213] && f[268]; // c9t609i60
	assign leaf[848] = f[709] && f[264] && f[213] && !f[712]; // c9t609i60
	assign leaf[849] = f[709] && f[264] && f[213] && f[712]; // c9t609i60
	assign leaf[850] = !f[740] && !f[462] && !f[457] && !f[181]; // c9t619i61
	assign leaf[851] = !f[740] && !f[462] && !f[457] && f[181]; // c9t619i61
	assign leaf[852] = !f[740] && !f[462] && f[457] && !f[375]; // c9t619i61
	assign leaf[853] = !f[740] && !f[462] && f[457] && f[375]; // c9t619i61
	assign leaf[854] = !f[740] && f[462] && !f[401] && !f[427]; // c9t619i61
	assign leaf[855] = !f[740] && f[462] && !f[401] && f[427]; // c9t619i61
	assign leaf[856] = !f[740] && f[462] && f[401] && !f[290]; // c9t619i61
	assign leaf[857] = !f[740] && f[462] && f[401] && f[290]; // c9t619i61
	assign leaf[858] = f[740] && !f[240] && !f[272]; // c9t619i61
	assign leaf[859] = f[740] && !f[240] && f[272]; // c9t619i61
	assign leaf[860] = f[740] && f[240] && !f[214] && !f[437]; // c9t619i61
	assign leaf[861] = f[740] && f[240] && !f[214] && f[437]; // c9t619i61
	assign leaf[862] = f[740] && f[240] && f[214] && !f[410]; // c9t619i61
	assign leaf[863] = f[740] && f[240] && f[214] && f[410]; // c9t619i61
	assign leaf[864] = !f[350] && !f[717] && !f[719] && !f[606]; // c9t629i62
	assign leaf[865] = !f[350] && !f[717] && !f[719] && f[606]; // c9t629i62
	assign leaf[866] = !f[350] && !f[717] && f[719] && !f[461]; // c9t629i62
	assign leaf[867] = !f[350] && !f[717] && f[719] && f[461]; // c9t629i62
	assign leaf[868] = !f[350] && f[717] && !f[237] && !f[608]; // c9t629i62
	assign leaf[869] = !f[350] && f[717] && !f[237] && f[608]; // c9t629i62
	assign leaf[870] = !f[350] && f[717] && f[237] && !f[378]; // c9t629i62
	assign leaf[871] = !f[350] && f[717] && f[237] && f[378]; // c9t629i62
	assign leaf[872] = f[350] && !f[488] && !f[324] && !f[373]; // c9t629i62
	assign leaf[873] = f[350] && !f[488] && !f[324] && f[373]; // c9t629i62
	assign leaf[874] = f[350] && !f[488] && f[324] && !f[187]; // c9t629i62
	assign leaf[875] = f[350] && !f[488] && f[324] && f[187]; // c9t629i62
	assign leaf[876] = f[350] && f[488] && !f[708] && !f[610]; // c9t629i62
	assign leaf[877] = f[350] && f[488] && !f[708] && f[610]; // c9t629i62
	assign leaf[878] = f[350] && f[488] && f[708] && !f[405]; // c9t629i62
	assign leaf[879] = f[350] && f[488] && f[708] && f[405]; // c9t629i62
	assign leaf[880] = !f[742] && !f[581] && !f[374] && !f[400]; // c9t639i63
	assign leaf[881] = !f[742] && !f[581] && !f[374] && f[400]; // c9t639i63
	assign leaf[882] = !f[742] && !f[581] && f[374] && !f[400]; // c9t639i63
	assign leaf[883] = !f[742] && !f[581] && f[374] && f[400]; // c9t639i63
	assign leaf[884] = !f[742] && f[581] && !f[496] && !f[580]; // c9t639i63
	assign leaf[885] = !f[742] && f[581] && !f[496] && f[580]; // c9t639i63
	assign leaf[886] = !f[742] && f[581] && f[496] && !f[411]; // c9t639i63
	assign leaf[887] = !f[742] && f[581] && f[496] && f[411]; // c9t639i63
	assign leaf[888] = f[742] && !f[326] && !f[319] && !f[406]; // c9t639i63
	assign leaf[889] = f[742] && !f[326] && !f[319] && f[406]; // c9t639i63
	assign leaf[890] = f[742] && !f[326] && f[319]; // c9t639i63
	assign leaf[891] = f[742] && f[326] && !f[351] && !f[487]; // c9t639i63
	assign leaf[892] = f[742] && f[326] && !f[351] && f[487]; // c9t639i63
	assign leaf[893] = f[742] && f[326] && f[351] && !f[660]; // c9t639i63
	assign leaf[894] = f[742] && f[326] && f[351] && f[660]; // c9t639i63
	assign leaf[895] = !f[717] && !f[718] && !f[128] && !f[517]; // c9t649i64
	assign leaf[896] = !f[717] && !f[718] && !f[128] && f[517]; // c9t649i64
	assign leaf[897] = !f[717] && !f[718] && f[128] && !f[575]; // c9t649i64
	assign leaf[898] = !f[717] && !f[718] && f[128] && f[575]; // c9t649i64
	assign leaf[899] = !f[717] && f[718] && !f[488] && !f[318]; // c9t649i64
	assign leaf[900] = !f[717] && f[718] && !f[488] && f[318]; // c9t649i64
	assign leaf[901] = !f[717] && f[718] && f[488] && !f[287]; // c9t649i64
	assign leaf[902] = !f[717] && f[718] && f[488] && f[287]; // c9t649i64
	assign leaf[903] = f[717] && !f[211] && !f[299] && !f[238]; // c9t649i64
	assign leaf[904] = f[717] && !f[211] && !f[299] && f[238]; // c9t649i64
	assign leaf[905] = f[717] && !f[211] && f[299] && !f[231]; // c9t649i64
	assign leaf[906] = f[717] && !f[211] && f[299] && f[231]; // c9t649i64
	assign leaf[907] = f[717] && f[211] && !f[691] && !f[212]; // c9t649i64
	assign leaf[908] = f[717] && f[211] && !f[691] && f[212]; // c9t649i64
	assign leaf[909] = f[717] && f[211] && f[691] && !f[438]; // c9t649i64
	assign leaf[910] = f[717] && f[211] && f[691] && f[438]; // c9t649i64
	assign leaf[911] = !f[687] && !f[509] && !f[584] && !f[320]; // c9t659i65
	assign leaf[912] = !f[687] && !f[509] && !f[584] && f[320]; // c9t659i65
	assign leaf[913] = !f[687] && !f[509] && f[584]; // c9t659i65
	assign leaf[914] = !f[687] && f[509] && !f[236]; // c9t659i65
	assign leaf[915] = !f[687] && f[509] && f[236] && !f[662]; // c9t659i65
	assign leaf[916] = !f[687] && f[509] && f[236] && f[662]; // c9t659i65
	assign leaf[917] = f[687] && !f[573] && !f[378] && !f[489]; // c9t659i65
	assign leaf[918] = f[687] && !f[573] && !f[378] && f[489]; // c9t659i65
	assign leaf[919] = f[687] && !f[573] && f[378] && !f[352]; // c9t659i65
	assign leaf[920] = f[687] && !f[573] && f[378] && f[352]; // c9t659i65
	assign leaf[921] = f[687] && f[573] && !f[158] && !f[484]; // c9t659i65
	assign leaf[922] = f[687] && f[573] && !f[158] && f[484]; // c9t659i65
	assign leaf[923] = f[687] && f[573] && f[158] && !f[428]; // c9t659i65
	assign leaf[924] = f[687] && f[573] && f[158] && f[428]; // c9t659i65
	assign leaf[925] = !f[368] && !f[498] && !f[184] && !f[240]; // c9t669i66
	assign leaf[926] = !f[368] && !f[498] && !f[184] && f[240]; // c9t669i66
	assign leaf[927] = !f[368] && !f[498] && f[184] && !f[240]; // c9t669i66
	assign leaf[928] = !f[368] && !f[498] && f[184] && f[240]; // c9t669i66
	assign leaf[929] = !f[368] && f[498] && !f[584] && !f[682]; // c9t669i66
	assign leaf[930] = !f[368] && f[498] && !f[584] && f[682]; // c9t669i66
	assign leaf[931] = !f[368] && f[498] && f[584]; // c9t669i66
	assign leaf[932] = f[368] && !f[347] && !f[385] && !f[520]; // c9t669i66
	assign leaf[933] = f[368] && !f[347] && !f[385] && f[520]; // c9t669i66
	assign leaf[934] = f[368] && !f[347] && f[385] && !f[398]; // c9t669i66
	assign leaf[935] = f[368] && !f[347] && f[385] && f[398]; // c9t669i66
	assign leaf[936] = f[368] && f[347] && !f[320]; // c9t669i66
	assign leaf[937] = f[368] && f[347] && f[320]; // c9t669i66
	assign leaf[938] = !f[351] && !f[383] && !f[381] && !f[519]; // c9t679i67
	assign leaf[939] = !f[351] && !f[383] && !f[381] && f[519]; // c9t679i67
	assign leaf[940] = !f[351] && !f[383] && f[381] && !f[270]; // c9t679i67
	assign leaf[941] = !f[351] && !f[383] && f[381] && f[270]; // c9t679i67
	assign leaf[942] = !f[351] && f[383] && !f[407] && !f[291]; // c9t679i67
	assign leaf[943] = !f[351] && f[383] && !f[407] && f[291]; // c9t679i67
	assign leaf[944] = !f[351] && f[383] && f[407] && !f[349]; // c9t679i67
	assign leaf[945] = !f[351] && f[383] && f[407] && f[349]; // c9t679i67
	assign leaf[946] = f[351] && !f[326] && !f[382] && !f[438]; // c9t679i67
	assign leaf[947] = f[351] && !f[326] && !f[382] && f[438]; // c9t679i67
	assign leaf[948] = f[351] && !f[326] && f[382] && !f[466]; // c9t679i67
	assign leaf[949] = f[351] && !f[326] && f[382] && f[466]; // c9t679i67
	assign leaf[950] = f[351] && f[326] && !f[213] && !f[600]; // c9t679i67
	assign leaf[951] = f[351] && f[326] && !f[213] && f[600]; // c9t679i67
	assign leaf[952] = f[351] && f[326] && f[213] && !f[538]; // c9t679i67
	assign leaf[953] = f[351] && f[326] && f[213] && f[538]; // c9t679i67
	assign leaf[954] = !f[323] && !f[401] && !f[427] && !f[375]; // c9t689i68
	assign leaf[955] = !f[323] && !f[401] && !f[427] && f[375]; // c9t689i68
	assign leaf[956] = !f[323] && !f[401] && f[427] && !f[497]; // c9t689i68
	assign leaf[957] = !f[323] && !f[401] && f[427] && f[497]; // c9t689i68
	assign leaf[958] = !f[323] && f[401] && !f[717] && !f[348]; // c9t689i68
	assign leaf[959] = !f[323] && f[401] && !f[717] && f[348]; // c9t689i68
	assign leaf[960] = !f[323] && f[401] && f[717] && !f[237]; // c9t689i68
	assign leaf[961] = !f[323] && f[401] && f[717] && f[237]; // c9t689i68
	assign leaf[962] = f[323] && !f[298] && !f[185] && !f[239]; // c9t689i68
	assign leaf[963] = f[323] && !f[298] && !f[185] && f[239]; // c9t689i68
	assign leaf[964] = f[323] && !f[298] && f[185] && !f[240]; // c9t689i68
	assign leaf[965] = f[323] && !f[298] && f[185] && f[240]; // c9t689i68
	assign leaf[966] = f[323] && f[298] && !f[245] && !f[209]; // c9t689i68
	assign leaf[967] = f[323] && f[298] && !f[245] && f[209]; // c9t689i68
	assign leaf[968] = f[323] && f[298] && f[245] && !f[405]; // c9t689i68
	assign leaf[969] = f[323] && f[298] && f[245] && f[405]; // c9t689i68
	assign leaf[970] = !f[500] && !f[350] && !f[438] && !f[522]; // c9t699i69
	assign leaf[971] = !f[500] && !f[350] && !f[438] && f[522]; // c9t699i69
	assign leaf[972] = !f[500] && !f[350] && f[438] && !f[493]; // c9t699i69
	assign leaf[973] = !f[500] && !f[350] && f[438] && f[493]; // c9t699i69
	assign leaf[974] = !f[500] && f[350] && !f[460] && !f[241]; // c9t699i69
	assign leaf[975] = !f[500] && f[350] && !f[460] && f[241]; // c9t699i69
	assign leaf[976] = !f[500] && f[350] && f[460] && !f[372]; // c9t699i69
	assign leaf[977] = !f[500] && f[350] && f[460] && f[372]; // c9t699i69
	assign leaf[978] = f[500]; // c9t699i69
	assign leaf[979] = !f[734] && !f[247] && !f[122] && !f[228]; // c9t709i70
	assign leaf[980] = !f[734] && !f[247] && !f[122] && f[228]; // c9t709i70
	assign leaf[981] = !f[734] && !f[247] && f[122]; // c9t709i70
	assign leaf[982] = !f[734] && f[247] && !f[215] && !f[514]; // c9t709i70
	assign leaf[983] = !f[734] && f[247] && !f[215] && f[514]; // c9t709i70
	assign leaf[984] = !f[734] && f[247] && f[215] && !f[404]; // c9t709i70
	assign leaf[985] = !f[734] && f[247] && f[215] && f[404]; // c9t709i70
	assign leaf[986] = f[734] && !f[624]; // c9t709i70
	assign leaf[987] = f[734] && f[624]; // c9t709i70
	assign leaf[988] = !f[566] && !f[175] && !f[639] && !f[524]; // c9t719i71
	assign leaf[989] = !f[566] && !f[175] && !f[639] && f[524]; // c9t719i71
	assign leaf[990] = !f[566] && !f[175] && f[639] && !f[426]; // c9t719i71
	assign leaf[991] = !f[566] && !f[175] && f[639] && f[426]; // c9t719i71
	assign leaf[992] = !f[566] && f[175] && !f[690]; // c9t719i71
	assign leaf[993] = !f[566] && f[175] && f[690]; // c9t719i71
	assign leaf[994] = f[566] && !f[551]; // c9t719i71
	assign leaf[995] = f[566] && f[551] && !f[320] && !f[315]; // c9t719i71
	assign leaf[996] = f[566] && f[551] && !f[320] && f[315]; // c9t719i71
	assign leaf[997] = f[566] && f[551] && f[320]; // c9t719i71
	assign leaf[998] = !f[381] && !f[432] && !f[491] && !f[206]; // c9t729i72
	assign leaf[999] = !f[381] && !f[432] && !f[491] && f[206]; // c9t729i72
	assign leaf[1000] = !f[381] && !f[432] && f[491] && !f[156]; // c9t729i72
	assign leaf[1001] = !f[381] && !f[432] && f[491] && f[156]; // c9t729i72
	assign leaf[1002] = !f[381] && f[432] && !f[374] && !f[460]; // c9t729i72
	assign leaf[1003] = !f[381] && f[432] && !f[374] && f[460]; // c9t729i72
	assign leaf[1004] = !f[381] && f[432] && f[374] && !f[514]; // c9t729i72
	assign leaf[1005] = !f[381] && f[432] && f[374] && f[514]; // c9t729i72
	assign leaf[1006] = f[381] && !f[437] && !f[520] && !f[263]; // c9t729i72
	assign leaf[1007] = f[381] && !f[437] && !f[520] && f[263]; // c9t729i72
	assign leaf[1008] = f[381] && !f[437] && f[520] && !f[490]; // c9t729i72
	assign leaf[1009] = f[381] && !f[437] && f[520] && f[490]; // c9t729i72
	assign leaf[1010] = f[381] && f[437] && !f[210] && !f[547]; // c9t729i72
	assign leaf[1011] = f[381] && f[437] && !f[210] && f[547]; // c9t729i72
	assign leaf[1012] = f[381] && f[437] && f[210] && !f[265]; // c9t729i72
	assign leaf[1013] = f[381] && f[437] && f[210] && f[265]; // c9t729i72
	assign leaf[1014] = !f[734] && !f[368] && !f[374] && !f[400]; // c9t739i73
	assign leaf[1015] = !f[734] && !f[368] && !f[374] && f[400]; // c9t739i73
	assign leaf[1016] = !f[734] && !f[368] && f[374] && !f[400]; // c9t739i73
	assign leaf[1017] = !f[734] && !f[368] && f[374] && f[400]; // c9t739i73
	assign leaf[1018] = !f[734] && f[368] && !f[347] && !f[270]; // c9t739i73
	assign leaf[1019] = !f[734] && f[368] && !f[347] && f[270]; // c9t739i73
	assign leaf[1020] = !f[734] && f[368] && f[347]; // c9t739i73
	assign leaf[1021] = f[734] && !f[321]; // c9t739i73
	assign leaf[1022] = f[734] && f[321]; // c9t739i73
	assign leaf[1023] = !f[351] && !f[377] && !f[323] && !f[407]; // c9t749i74
	assign leaf[1024] = !f[351] && !f[377] && !f[323] && f[407]; // c9t749i74
	assign leaf[1025] = !f[351] && !f[377] && f[323] && !f[709]; // c9t749i74
	assign leaf[1026] = !f[351] && !f[377] && f[323] && f[709]; // c9t749i74
	assign leaf[1027] = !f[351] && f[377] && !f[652] && !f[713]; // c9t749i74
	assign leaf[1028] = !f[351] && f[377] && !f[652] && f[713]; // c9t749i74
	assign leaf[1029] = !f[351] && f[377] && f[652] && !f[412]; // c9t749i74
	assign leaf[1030] = !f[351] && f[377] && f[652] && f[412]; // c9t749i74
	assign leaf[1031] = f[351] && !f[511] && !f[434] && !f[152]; // c9t749i74
	assign leaf[1032] = f[351] && !f[511] && !f[434] && f[152]; // c9t749i74
	assign leaf[1033] = f[351] && !f[511] && f[434] && !f[320]; // c9t749i74
	assign leaf[1034] = f[351] && !f[511] && f[434] && f[320]; // c9t749i74
	assign leaf[1035] = f[351] && f[511] && !f[659] && !f[260]; // c9t749i74
	assign leaf[1036] = f[351] && f[511] && !f[659] && f[260]; // c9t749i74
	assign leaf[1037] = f[351] && f[511] && f[659] && !f[521]; // c9t749i74
	assign leaf[1038] = f[351] && f[511] && f[659] && f[521]; // c9t749i74
	assign leaf[1039] = !f[686] && !f[603] && !f[715] && !f[186]; // c9t759i75
	assign leaf[1040] = !f[686] && !f[603] && !f[715] && f[186]; // c9t759i75
	assign leaf[1041] = !f[686] && !f[603] && f[715] && !f[521]; // c9t759i75
	assign leaf[1042] = !f[686] && !f[603] && f[715] && f[521]; // c9t759i75
	assign leaf[1043] = !f[686] && f[603] && !f[181] && !f[744]; // c9t759i75
	assign leaf[1044] = !f[686] && f[603] && !f[181] && f[744]; // c9t759i75
	assign leaf[1045] = !f[686] && f[603] && f[181] && !f[659]; // c9t759i75
	assign leaf[1046] = !f[686] && f[603] && f[181] && f[659]; // c9t759i75
	assign leaf[1047] = f[686] && !f[572] && !f[518] && !f[547]; // c9t759i75
	assign leaf[1048] = f[686] && !f[572] && !f[518] && f[547]; // c9t759i75
	assign leaf[1049] = f[686] && !f[572] && f[518] && !f[264]; // c9t759i75
	assign leaf[1050] = f[686] && !f[572] && f[518] && f[264]; // c9t759i75
	assign leaf[1051] = f[686] && f[572] && !f[428] && !f[489]; // c9t759i75
	assign leaf[1052] = f[686] && f[572] && !f[428] && f[489]; // c9t759i75
	assign leaf[1053] = f[686] && f[572] && f[428] && !f[604]; // c9t759i75
	assign leaf[1054] = f[686] && f[572] && f[428] && f[604]; // c9t759i75
	assign leaf[1055] = !f[742] && !f[162] && !f[229] && !f[740]; // c9t769i76
	assign leaf[1056] = !f[742] && !f[162] && !f[229] && f[740]; // c9t769i76
	assign leaf[1057] = !f[742] && !f[162] && f[229] && !f[260]; // c9t769i76
	assign leaf[1058] = !f[742] && !f[162] && f[229] && f[260]; // c9t769i76
	assign leaf[1059] = !f[742] && f[162] && !f[246]; // c9t769i76
	assign leaf[1060] = !f[742] && f[162] && f[246]; // c9t769i76
	assign leaf[1061] = f[742] && !f[328] && !f[259] && !f[326]; // c9t769i76
	assign leaf[1062] = f[742] && !f[328] && !f[259] && f[326]; // c9t769i76
	assign leaf[1063] = f[742] && !f[328] && f[259]; // c9t769i76
	assign leaf[1064] = f[742] && f[328] && !f[345]; // c9t769i76
	assign leaf[1065] = f[742] && f[328] && f[345] && !f[494]; // c9t769i76
	assign leaf[1066] = f[742] && f[328] && f[345] && f[494]; // c9t769i76
	assign leaf[1067] = !f[350] && !f[384] && !f[467] && !f[378]; // c9t779i77
	assign leaf[1068] = !f[350] && !f[384] && !f[467] && f[378]; // c9t779i77
	assign leaf[1069] = !f[350] && !f[384] && f[467] && !f[288]; // c9t779i77
	assign leaf[1070] = !f[350] && !f[384] && f[467] && f[288]; // c9t779i77
	assign leaf[1071] = !f[350] && f[384] && !f[467] && !f[215]; // c9t779i77
	assign leaf[1072] = !f[350] && f[384] && !f[467] && f[215]; // c9t779i77
	assign leaf[1073] = !f[350] && f[384] && f[467] && !f[246]; // c9t779i77
	assign leaf[1074] = !f[350] && f[384] && f[467] && f[246]; // c9t779i77
	assign leaf[1075] = f[350] && !f[324] && !f[651] && !f[352]; // c9t779i77
	assign leaf[1076] = f[350] && !f[324] && !f[651] && f[352]; // c9t779i77
	assign leaf[1077] = f[350] && !f[324] && f[651]; // c9t779i77
	assign leaf[1078] = f[350] && f[324] && !f[487] && !f[384]; // c9t779i77
	assign leaf[1079] = f[350] && f[324] && !f[487] && f[384]; // c9t779i77
	assign leaf[1080] = f[350] && f[324] && f[487] && !f[628]; // c9t779i77
	assign leaf[1081] = f[350] && f[324] && f[487] && f[628]; // c9t779i77
	assign leaf[1082] = !f[575] && !f[294] && !f[685] && !f[345]; // c9t789i78
	assign leaf[1083] = !f[575] && !f[294] && !f[685] && f[345]; // c9t789i78
	assign leaf[1084] = !f[575] && !f[294] && f[685] && !f[520]; // c9t789i78
	assign leaf[1085] = !f[575] && !f[294] && f[685] && f[520]; // c9t789i78
	assign leaf[1086] = !f[575] && f[294] && !f[301] && !f[259]; // c9t789i78
	assign leaf[1087] = !f[575] && f[294] && !f[301] && f[259]; // c9t789i78
	assign leaf[1088] = !f[575] && f[294] && f[301] && !f[433]; // c9t789i78
	assign leaf[1089] = !f[575] && f[294] && f[301] && f[433]; // c9t789i78
	assign leaf[1090] = f[575] && !f[517] && !f[209] && !f[181]; // c9t789i78
	assign leaf[1091] = f[575] && !f[517] && !f[209] && f[181]; // c9t789i78
	assign leaf[1092] = f[575] && !f[517] && f[209] && !f[456]; // c9t789i78
	assign leaf[1093] = f[575] && !f[517] && f[209] && f[456]; // c9t789i78
	assign leaf[1094] = f[575] && f[517] && !f[456] && !f[458]; // c9t789i78
	assign leaf[1095] = f[575] && f[517] && !f[456] && f[458]; // c9t789i78
	assign leaf[1096] = f[575] && f[517] && f[456] && !f[657]; // c9t789i78
	assign leaf[1097] = f[575] && f[517] && f[456] && f[657]; // c9t789i78
	assign leaf[1098] = !f[131] && !f[599] && !f[377] && !f[488]; // c9t799i79
	assign leaf[1099] = !f[131] && !f[599] && !f[377] && f[488]; // c9t799i79
	assign leaf[1100] = !f[131] && !f[599] && f[377] && !f[714]; // c9t799i79
	assign leaf[1101] = !f[131] && !f[599] && f[377] && f[714]; // c9t799i79
	assign leaf[1102] = !f[131] && f[599] && !f[487] && !f[378]; // c9t799i79
	assign leaf[1103] = !f[131] && f[599] && !f[487] && f[378]; // c9t799i79
	assign leaf[1104] = !f[131] && f[599] && f[487] && !f[434]; // c9t799i79
	assign leaf[1105] = !f[131] && f[599] && f[487] && f[434]; // c9t799i79
	assign leaf[1106] = f[131]; // c9t799i79
	assign leaf[1107] = !f[244] && !f[275] && !f[327] && !f[213]; // c9t809i80
	assign leaf[1108] = !f[244] && !f[275] && !f[327] && f[213]; // c9t809i80
	assign leaf[1109] = !f[244] && !f[275] && f[327] && !f[211]; // c9t809i80
	assign leaf[1110] = !f[244] && !f[275] && f[327] && f[211]; // c9t809i80
	assign leaf[1111] = !f[244] && f[275] && !f[214]; // c9t809i80
	assign leaf[1112] = !f[244] && f[275] && f[214]; // c9t809i80
	assign leaf[1113] = f[244] && !f[385] && !f[209] && !f[299]; // c9t809i80
	assign leaf[1114] = f[244] && !f[385] && !f[209] && f[299]; // c9t809i80
	assign leaf[1115] = f[244] && !f[385] && f[209] && !f[185]; // c9t809i80
	assign leaf[1116] = f[244] && !f[385] && f[209] && f[185]; // c9t809i80
	assign leaf[1117] = f[244] && f[385] && !f[440] && !f[274]; // c9t809i80
	assign leaf[1118] = f[244] && f[385] && !f[440] && f[274]; // c9t809i80
	assign leaf[1119] = f[244] && f[385] && f[440] && !f[486]; // c9t809i80
	assign leaf[1120] = f[244] && f[385] && f[440] && f[486]; // c9t809i80
	assign leaf[1121] = !f[201] && !f[632] && !f[128] && !f[292]; // c9t819i81
	assign leaf[1122] = !f[201] && !f[632] && !f[128] && f[292]; // c9t819i81
	assign leaf[1123] = !f[201] && !f[632] && f[128]; // c9t819i81
	assign leaf[1124] = !f[201] && f[632] && !f[546] && !f[155]; // c9t819i81
	assign leaf[1125] = !f[201] && f[632] && !f[546] && f[155]; // c9t819i81
	assign leaf[1126] = !f[201] && f[632] && f[546] && !f[513]; // c9t819i81
	assign leaf[1127] = !f[201] && f[632] && f[546] && f[513]; // c9t819i81
	assign leaf[1128] = f[201] && !f[428]; // c9t819i81
	assign leaf[1129] = f[201] && f[428]; // c9t819i81
	assign leaf[1130] = !f[599] && !f[543] && !f[540] && !f[740]; // c9t829i82
	assign leaf[1131] = !f[599] && !f[543] && !f[540] && f[740]; // c9t829i82
	assign leaf[1132] = !f[599] && !f[543] && f[540] && !f[482]; // c9t829i82
	assign leaf[1133] = !f[599] && !f[543] && f[540] && f[482]; // c9t829i82
	assign leaf[1134] = !f[599] && f[543] && !f[432] && !f[459]; // c9t829i82
	assign leaf[1135] = !f[599] && f[543] && !f[432] && f[459]; // c9t829i82
	assign leaf[1136] = !f[599] && f[543] && f[432] && !f[428]; // c9t829i82
	assign leaf[1137] = !f[599] && f[543] && f[432] && f[428]; // c9t829i82
	assign leaf[1138] = f[599] && !f[488] && !f[272] && !f[511]; // c9t829i82
	assign leaf[1139] = f[599] && !f[488] && !f[272] && f[511]; // c9t829i82
	assign leaf[1140] = f[599] && !f[488] && f[272] && !f[238]; // c9t829i82
	assign leaf[1141] = f[599] && !f[488] && f[272] && f[238]; // c9t829i82
	assign leaf[1142] = f[599] && f[488] && !f[186] && !f[516]; // c9t829i82
	assign leaf[1143] = f[599] && f[488] && !f[186] && f[516]; // c9t829i82
	assign leaf[1144] = f[599] && f[488] && f[186] && !f[680]; // c9t829i82
	assign leaf[1145] = f[599] && f[488] && f[186] && f[680]; // c9t829i82
	assign leaf[1146] = !f[744] && !f[524] && !f[469] && !f[379]; // c9t839i83
	assign leaf[1147] = !f[744] && !f[524] && !f[469] && f[379]; // c9t839i83
	assign leaf[1148] = !f[744] && !f[524] && f[469] && !f[413]; // c9t839i83
	assign leaf[1149] = !f[744] && !f[524] && f[469] && f[413]; // c9t839i83
	assign leaf[1150] = !f[744] && f[524] && !f[259] && !f[565]; // c9t839i83
	assign leaf[1151] = !f[744] && f[524] && !f[259] && f[565]; // c9t839i83
	assign leaf[1152] = !f[744] && f[524] && f[259] && !f[290]; // c9t839i83
	assign leaf[1153] = !f[744] && f[524] && f[259] && f[290]; // c9t839i83
	assign leaf[1154] = f[744] && !f[434] && !f[322] && !f[351]; // c9t839i83
	assign leaf[1155] = f[744] && !f[434] && !f[322] && f[351]; // c9t839i83
	assign leaf[1156] = f[744] && !f[434] && f[322]; // c9t839i83
	assign leaf[1157] = f[744] && f[434] && !f[690] && !f[287]; // c9t839i83
	assign leaf[1158] = f[744] && f[434] && !f[690] && f[287]; // c9t839i83
	assign leaf[1159] = f[744] && f[434] && f[690]; // c9t839i83
	assign leaf[1160] = !f[508] && !f[350] && !f[340] && !f[401]; // c9t849i84
	assign leaf[1161] = !f[508] && !f[350] && !f[340] && f[401]; // c9t849i84
	assign leaf[1162] = !f[508] && !f[350] && f[340] && !f[212]; // c9t849i84
	assign leaf[1163] = !f[508] && !f[350] && f[340] && f[212]; // c9t849i84
	assign leaf[1164] = !f[508] && f[350] && !f[352] && !f[267]; // c9t849i84
	assign leaf[1165] = !f[508] && f[350] && !f[352] && f[267]; // c9t849i84
	assign leaf[1166] = !f[508] && f[350] && f[352] && !f[402]; // c9t849i84
	assign leaf[1167] = !f[508] && f[350] && f[352] && f[402]; // c9t849i84
	assign leaf[1168] = f[508]; // c9t849i84
	assign leaf[1169] = !f[742] && !f[407] && !f[346] && !f[574]; // c9t859i85
	assign leaf[1170] = !f[742] && !f[407] && !f[346] && f[574]; // c9t859i85
	assign leaf[1171] = !f[742] && !f[407] && f[346] && !f[432]; // c9t859i85
	assign leaf[1172] = !f[742] && !f[407] && f[346] && f[432]; // c9t859i85
	assign leaf[1173] = !f[742] && f[407] && !f[291] && !f[211]; // c9t859i85
	assign leaf[1174] = !f[742] && f[407] && !f[291] && f[211]; // c9t859i85
	assign leaf[1175] = !f[742] && f[407] && f[291] && !f[206]; // c9t859i85
	assign leaf[1176] = !f[742] && f[407] && f[291] && f[206]; // c9t859i85
	assign leaf[1177] = f[742] && !f[573] && !f[315] && !f[379]; // c9t859i85
	assign leaf[1178] = f[742] && !f[573] && !f[315] && f[379]; // c9t859i85
	assign leaf[1179] = f[742] && !f[573] && f[315] && !f[209]; // c9t859i85
	assign leaf[1180] = f[742] && !f[573] && f[315] && f[209]; // c9t859i85
	assign leaf[1181] = f[742] && f[573] && !f[458]; // c9t859i85
	assign leaf[1182] = f[742] && f[573] && f[458]; // c9t859i85
	assign leaf[1183] = !f[500] && !f[162] && !f[122] && !f[686]; // c9t869i86
	assign leaf[1184] = !f[500] && !f[162] && !f[122] && f[686]; // c9t869i86
	assign leaf[1185] = !f[500] && !f[162] && f[122]; // c9t869i86
	assign leaf[1186] = !f[500] && f[162]; // c9t869i86
	assign leaf[1187] = f[500]; // c9t869i86
	assign leaf[1188] = !f[742] && !f[351] && !f[433] && !f[489]; // c9t879i87
	assign leaf[1189] = !f[742] && !f[351] && !f[433] && f[489]; // c9t879i87
	assign leaf[1190] = !f[742] && !f[351] && f[433] && !f[516]; // c9t879i87
	assign leaf[1191] = !f[742] && !f[351] && f[433] && f[516]; // c9t879i87
	assign leaf[1192] = !f[742] && f[351] && !f[353] && !f[409]; // c9t879i87
	assign leaf[1193] = !f[742] && f[351] && !f[353] && f[409]; // c9t879i87
	assign leaf[1194] = !f[742] && f[351] && f[353] && !f[385]; // c9t879i87
	assign leaf[1195] = !f[742] && f[351] && f[353] && f[385]; // c9t879i87
	assign leaf[1196] = f[742] && !f[290] && !f[407]; // c9t879i87
	assign leaf[1197] = f[742] && !f[290] && f[407] && !f[294]; // c9t879i87
	assign leaf[1198] = f[742] && !f[290] && f[407] && f[294]; // c9t879i87
	assign leaf[1199] = f[742] && f[290] && !f[234] && !f[399]; // c9t879i87
	assign leaf[1200] = f[742] && f[290] && !f[234] && f[399]; // c9t879i87
	assign leaf[1201] = f[742] && f[290] && f[234] && !f[461]; // c9t879i87
	assign leaf[1202] = f[742] && f[290] && f[234] && f[461]; // c9t879i87
	assign leaf[1203] = !f[269] && !f[185] && !f[299] && !f[412]; // c9t889i88
	assign leaf[1204] = !f[269] && !f[185] && !f[299] && f[412]; // c9t889i88
	assign leaf[1205] = !f[269] && !f[185] && f[299] && !f[241]; // c9t889i88
	assign leaf[1206] = !f[269] && !f[185] && f[299] && f[241]; // c9t889i88
	assign leaf[1207] = !f[269] && f[185] && !f[212] && !f[657]; // c9t889i88
	assign leaf[1208] = !f[269] && f[185] && !f[212] && f[657]; // c9t889i88
	assign leaf[1209] = !f[269] && f[185] && f[212] && !f[156]; // c9t889i88
	assign leaf[1210] = !f[269] && f[185] && f[212] && f[156]; // c9t889i88
	assign leaf[1211] = f[269] && !f[187] && !f[322] && !f[486]; // c9t889i88
	assign leaf[1212] = f[269] && !f[187] && !f[322] && f[486]; // c9t889i88
	assign leaf[1213] = f[269] && !f[187] && f[322] && !f[403]; // c9t889i88
	assign leaf[1214] = f[269] && !f[187] && f[322] && f[403]; // c9t889i88
	assign leaf[1215] = f[269] && f[187] && !f[185] && !f[540]; // c9t889i88
	assign leaf[1216] = f[269] && f[187] && !f[185] && f[540]; // c9t889i88
	assign leaf[1217] = f[269] && f[187] && f[185] && !f[241]; // c9t889i88
	assign leaf[1218] = f[269] && f[187] && f[185] && f[241]; // c9t889i88
	assign leaf[1219] = !f[183] && !f[239] && !f[657] && !f[291]; // c9t899i89
	assign leaf[1220] = !f[183] && !f[239] && !f[657] && f[291]; // c9t899i89
	assign leaf[1221] = !f[183] && !f[239] && f[657] && !f[156]; // c9t899i89
	assign leaf[1222] = !f[183] && !f[239] && f[657] && f[156]; // c9t899i89
	assign leaf[1223] = !f[183] && f[239] && !f[433] && !f[381]; // c9t899i89
	assign leaf[1224] = !f[183] && f[239] && !f[433] && f[381]; // c9t899i89
	assign leaf[1225] = !f[183] && f[239] && f[433] && !f[462]; // c9t899i89
	assign leaf[1226] = !f[183] && f[239] && f[433] && f[462]; // c9t899i89
	assign leaf[1227] = f[183] && !f[211] && !f[398] && !f[184]; // c9t899i89
	assign leaf[1228] = f[183] && !f[211] && !f[398] && f[184]; // c9t899i89
	assign leaf[1229] = f[183] && !f[211] && f[398]; // c9t899i89
	assign leaf[1230] = f[183] && f[211] && !f[291] && !f[206]; // c9t899i89
	assign leaf[1231] = f[183] && f[211] && !f[291] && f[206]; // c9t899i89
	assign leaf[1232] = f[183] && f[211] && f[291] && !f[345]; // c9t899i89
	assign leaf[1233] = f[183] && f[211] && f[291] && f[345]; // c9t899i89
	assign leaf[1234] = !f[256] && !f[342] && !f[387] && !f[320]; // c9t909i90
	assign leaf[1235] = !f[256] && !f[342] && !f[387] && f[320]; // c9t909i90
	assign leaf[1236] = !f[256] && !f[342] && f[387]; // c9t909i90
	assign leaf[1237] = !f[256] && f[342] && !f[290] && !f[687]; // c9t909i90
	assign leaf[1238] = !f[256] && f[342] && !f[290] && f[687]; // c9t909i90
	assign leaf[1239] = !f[256] && f[342] && f[290] && !f[454]; // c9t909i90
	assign leaf[1240] = !f[256] && f[342] && f[290] && f[454]; // c9t909i90
	assign leaf[1241] = f[256] && !f[398]; // c9t909i90
	assign leaf[1242] = f[256] && f[398]; // c9t909i90
	assign leaf[1243] = !f[742] && !f[740] && !f[182] && !f[266]; // c9t919i91
	assign leaf[1244] = !f[742] && !f[740] && !f[182] && f[266]; // c9t919i91
	assign leaf[1245] = !f[742] && !f[740] && f[182] && !f[237]; // c9t919i91
	assign leaf[1246] = !f[742] && !f[740] && f[182] && f[237]; // c9t919i91
	assign leaf[1247] = !f[742] && f[740] && !f[406] && !f[461]; // c9t919i91
	assign leaf[1248] = !f[742] && f[740] && !f[406] && f[461]; // c9t919i91
	assign leaf[1249] = !f[742] && f[740] && f[406] && !f[289]; // c9t919i91
	assign leaf[1250] = !f[742] && f[740] && f[406] && f[289]; // c9t919i91
	assign leaf[1251] = f[742] && !f[326] && !f[319]; // c9t919i91
	assign leaf[1252] = f[742] && !f[326] && f[319]; // c9t919i91
	assign leaf[1253] = f[742] && f[326] && !f[601] && !f[458]; // c9t919i91
	assign leaf[1254] = f[742] && f[326] && !f[601] && f[458]; // c9t919i91
	assign leaf[1255] = f[742] && f[326] && f[601]; // c9t919i91
	assign leaf[1256] = !f[740] && !f[472] && !f[184] && !f[602]; // c9t929i92
	assign leaf[1257] = !f[740] && !f[472] && !f[184] && f[602]; // c9t929i92
	assign leaf[1258] = !f[740] && !f[472] && f[184] && !f[717]; // c9t929i92
	assign leaf[1259] = !f[740] && !f[472] && f[184] && f[717]; // c9t929i92
	assign leaf[1260] = !f[740] && f[472]; // c9t929i92
	assign leaf[1261] = f[740] && !f[544] && !f[490] && !f[290]; // c9t929i92
	assign leaf[1262] = f[740] && !f[544] && !f[490] && f[290]; // c9t929i92
	assign leaf[1263] = f[740] && !f[544] && f[490] && !f[713]; // c9t929i92
	assign leaf[1264] = f[740] && !f[544] && f[490] && f[713]; // c9t929i92
	assign leaf[1265] = f[740] && f[544]; // c9t929i92
	assign leaf[1266] = !f[201] && !f[575] && !f[685] && !f[349]; // c9t939i93
	assign leaf[1267] = !f[201] && !f[575] && !f[685] && f[349]; // c9t939i93
	assign leaf[1268] = !f[201] && !f[575] && f[685] && !f[294]; // c9t939i93
	assign leaf[1269] = !f[201] && !f[575] && f[685] && f[294]; // c9t939i93
	assign leaf[1270] = !f[201] && f[575] && !f[518] && !f[459]; // c9t939i93
	assign leaf[1271] = !f[201] && f[575] && !f[518] && f[459]; // c9t939i93
	assign leaf[1272] = !f[201] && f[575] && f[518] && !f[179]; // c9t939i93
	assign leaf[1273] = !f[201] && f[575] && f[518] && f[179]; // c9t939i93
	assign leaf[1274] = f[201]; // c9t939i93
	assign leaf[1275] = !f[536] && !f[201] && !f[599] && !f[654]; // c9t949i94
	assign leaf[1276] = !f[536] && !f[201] && !f[599] && f[654]; // c9t949i94
	assign leaf[1277] = !f[536] && !f[201] && f[599] && !f[487]; // c9t949i94
	assign leaf[1278] = !f[536] && !f[201] && f[599] && f[487]; // c9t949i94
	assign leaf[1279] = !f[536] && f[201]; // c9t949i94
	assign leaf[1280] = f[536]; // c9t949i94
	assign leaf[1281] = !f[174] && !f[322] && !f[402] && !f[456]; // c9t959i95
	assign leaf[1282] = !f[174] && !f[322] && !f[402] && f[456]; // c9t959i95
	assign leaf[1283] = !f[174] && !f[322] && f[402] && !f[455]; // c9t959i95
	assign leaf[1284] = !f[174] && !f[322] && f[402] && f[455]; // c9t959i95
	assign leaf[1285] = !f[174] && f[322] && !f[157] && !f[540]; // c9t959i95
	assign leaf[1286] = !f[174] && f[322] && !f[157] && f[540]; // c9t959i95
	assign leaf[1287] = !f[174] && f[322] && f[157] && !f[315]; // c9t959i95
	assign leaf[1288] = !f[174] && f[322] && f[157] && f[315]; // c9t959i95
	assign leaf[1289] = f[174]; // c9t959i95
	assign leaf[1290] = !f[408] && !f[468] && !f[157] && !f[410]; // c9t969i96
	assign leaf[1291] = !f[408] && !f[468] && !f[157] && f[410]; // c9t969i96
	assign leaf[1292] = !f[408] && !f[468] && f[157] && !f[521]; // c9t969i96
	assign leaf[1293] = !f[408] && !f[468] && f[157] && f[521]; // c9t969i96
	assign leaf[1294] = !f[408] && f[468] && !f[517] && !f[574]; // c9t969i96
	assign leaf[1295] = !f[408] && f[468] && !f[517] && f[574]; // c9t969i96
	assign leaf[1296] = !f[408] && f[468] && f[517] && !f[470]; // c9t969i96
	assign leaf[1297] = !f[408] && f[468] && f[517] && f[470]; // c9t969i96
	assign leaf[1298] = f[408] && !f[467] && !f[412] && !f[352]; // c9t969i96
	assign leaf[1299] = f[408] && !f[467] && !f[412] && f[352]; // c9t969i96
	assign leaf[1300] = f[408] && !f[467] && f[412] && !f[328]; // c9t969i96
	assign leaf[1301] = f[408] && !f[467] && f[412] && f[328]; // c9t969i96
	assign leaf[1302] = f[408] && f[467] && !f[384] && !f[635]; // c9t969i96
	assign leaf[1303] = f[408] && f[467] && !f[384] && f[635]; // c9t969i96
	assign leaf[1304] = f[408] && f[467] && f[384] && !f[322]; // c9t969i96
	assign leaf[1305] = f[408] && f[467] && f[384] && f[322]; // c9t969i96
	assign leaf[1306] = !f[191] && !f[326] && !f[396] && !f[462]; // c9t979i97
	assign leaf[1307] = !f[191] && !f[326] && !f[396] && f[462]; // c9t979i97
	assign leaf[1308] = !f[191] && !f[326] && f[396] && !f[398]; // c9t979i97
	assign leaf[1309] = !f[191] && !f[326] && f[396] && f[398]; // c9t979i97
	assign leaf[1310] = !f[191] && f[326] && !f[271] && !f[330]; // c9t979i97
	assign leaf[1311] = !f[191] && f[326] && !f[271] && f[330]; // c9t979i97
	assign leaf[1312] = !f[191] && f[326] && f[271] && !f[356]; // c9t979i97
	assign leaf[1313] = !f[191] && f[326] && f[271] && f[356]; // c9t979i97
	assign leaf[1314] = f[191] && !f[188]; // c9t979i97
	assign leaf[1315] = f[191] && f[188]; // c9t979i97
	assign leaf[1316] = !f[186] && !f[262] && !f[205] && !f[466]; // c9t989i98
	assign leaf[1317] = !f[186] && !f[262] && !f[205] && f[466]; // c9t989i98
	assign leaf[1318] = !f[186] && !f[262] && f[205] && !f[179]; // c9t989i98
	assign leaf[1319] = !f[186] && !f[262] && f[205] && f[179]; // c9t989i98
	assign leaf[1320] = !f[186] && f[262] && !f[246] && !f[235]; // c9t989i98
	assign leaf[1321] = !f[186] && f[262] && !f[246] && f[235]; // c9t989i98
	assign leaf[1322] = !f[186] && f[262] && f[246] && !f[207]; // c9t989i98
	assign leaf[1323] = !f[186] && f[262] && f[246] && f[207]; // c9t989i98
	assign leaf[1324] = f[186] && !f[241] && !f[185] && !f[263]; // c9t989i98
	assign leaf[1325] = f[186] && !f[241] && !f[185] && f[263]; // c9t989i98
	assign leaf[1326] = f[186] && !f[241] && f[185] && !f[684]; // c9t989i98
	assign leaf[1327] = f[186] && !f[241] && f[185] && f[684]; // c9t989i98
	assign leaf[1328] = f[186] && f[241] && !f[238] && !f[183]; // c9t989i98
	assign leaf[1329] = f[186] && f[241] && !f[238] && f[183]; // c9t989i98
	assign leaf[1330] = f[186] && f[241] && f[238] && !f[491]; // c9t989i98
	assign leaf[1331] = f[186] && f[241] && f[238] && f[491]; // c9t989i98
	assign leaf[1332] = !f[350] && !f[322] && !f[410] && !f[206]; // c9t999i99
	assign leaf[1333] = !f[350] && !f[322] && !f[410] && f[206]; // c9t999i99
	assign leaf[1334] = !f[350] && !f[322] && f[410] && !f[407]; // c9t999i99
	assign leaf[1335] = !f[350] && !f[322] && f[410] && f[407]; // c9t999i99
	assign leaf[1336] = !f[350] && f[322] && !f[266] && !f[352]; // c9t999i99
	assign leaf[1337] = !f[350] && f[322] && !f[266] && f[352]; // c9t999i99
	assign leaf[1338] = !f[350] && f[322] && f[266] && !f[238]; // c9t999i99
	assign leaf[1339] = !f[350] && f[322] && f[266] && f[238]; // c9t999i99
	assign leaf[1340] = f[350] && !f[324] && !f[430] && !f[204]; // c9t999i99
	assign leaf[1341] = f[350] && !f[324] && !f[430] && f[204]; // c9t999i99
	assign leaf[1342] = f[350] && !f[324] && f[430] && !f[211]; // c9t999i99
	assign leaf[1343] = f[350] && !f[324] && f[430] && f[211]; // c9t999i99
	assign leaf[1344] = f[350] && f[324] && !f[237] && !f[180]; // c9t999i99
	assign leaf[1345] = f[350] && f[324] && !f[237] && f[180]; // c9t999i99
	assign leaf[1346] = f[350] && f[324] && f[237] && !f[180]; // c9t999i99
	assign leaf[1347] = f[350] && f[324] && f[237] && f[180]; // c9t999i99
endmodule