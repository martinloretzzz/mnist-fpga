module decision_tree_leaves(input logic [0:783] f, output logic [0:13595] leaf);
// Tree 0, Classifier 0, Iteration: 0
	assign leaf[0] = !f[358] && !f[357] && !f[359] && !f[384];
	assign leaf[1] = !f[358] && !f[357] && !f[359] && f[384];
	assign leaf[2] = !f[358] && !f[357] && f[359] && !f[462];
	assign leaf[3] = !f[358] && !f[357] && f[359] && f[462];
	assign leaf[4] = !f[358] && f[357] && !f[435] && !f[512];
	assign leaf[5] = !f[358] && f[357] && !f[435] && f[512];
	assign leaf[6] = !f[358] && f[357] && f[435] && !f[322];
	assign leaf[7] = !f[358] && f[357] && f[435] && f[322];
	assign leaf[8] = f[358] && !f[435] && !f[596] && !f[213];
	assign leaf[9] = f[358] && !f[435] && !f[596] && f[213];
	assign leaf[10] = f[358] && !f[435] && f[596] && !f[461];
	assign leaf[11] = f[358] && !f[435] && f[596] && f[461];
	assign leaf[12] = f[358] && f[435] && !f[295] && !f[245];
	assign leaf[13] = f[358] && f[435] && !f[295] && f[245];
	assign leaf[14] = f[358] && f[435] && f[295] && !f[538];
	assign leaf[15] = f[358] && f[435] && f[295] && f[538];
	
	// Tree 1, Classifier 1, Iteration: 0
	assign leaf[16] = !f[350] && !f[351] && !f[349];
	assign leaf[17] = !f[350] && !f[351] && f[349] && !f[347];
	assign leaf[18] = !f[350] && !f[351] && f[349] && f[347];
	assign leaf[19] = !f[350] && f[351] && !f[236] && !f[492];
	assign leaf[20] = !f[350] && f[351] && !f[236] && f[492];
	assign leaf[21] = !f[350] && f[351] && f[236] && !f[608];
	assign leaf[22] = !f[350] && f[351] && f[236] && f[608];
	assign leaf[23] = f[350] && !f[489] && !f[490] && !f[488];
	assign leaf[24] = f[350] && !f[489] && !f[490] && f[488];
	assign leaf[25] = f[350] && !f[489] && f[490] && !f[404];
	assign leaf[26] = f[350] && !f[489] && f[490] && f[404];
	assign leaf[27] = f[350] && f[489] && !f[521] && !f[375];
	assign leaf[28] = f[350] && f[489] && !f[521] && f[375];
	assign leaf[29] = f[350] && f[489] && f[521] && !f[487];
	assign leaf[30] = f[350] && f[489] && f[521] && f[487];
	
	// Tree 2, Classifier 2, Iteration: 0
	assign leaf[31] = !f[583] && !f[124] && !f[528] && !f[564];
	assign leaf[32] = !f[583] && !f[124] && !f[528] && f[564];
	assign leaf[33] = !f[583] && !f[124] && f[528] && !f[371];
	assign leaf[34] = !f[583] && !f[124] && f[528] && f[371];
	assign leaf[35] = !f[583] && f[124] && !f[346] && !f[349];
	assign leaf[36] = !f[583] && f[124] && !f[346] && f[349];
	assign leaf[37] = !f[583] && f[124] && f[346] && !f[93];
	assign leaf[38] = !f[583] && f[124] && f[346] && f[93];
	assign leaf[39] = f[583] && !f[343] && !f[346] && !f[369];
	assign leaf[40] = f[583] && !f[343] && !f[346] && f[369];
	assign leaf[41] = f[583] && !f[343] && f[346] && !f[520];
	assign leaf[42] = f[583] && !f[343] && f[346] && f[520];
	assign leaf[43] = f[583] && f[343] && !f[519] && !f[517];
	assign leaf[44] = f[583] && f[343] && !f[519] && f[517];
	assign leaf[45] = f[583] && f[343] && f[519] && !f[442];
	assign leaf[46] = f[583] && f[343] && f[519] && f[442];
	
	// Tree 3, Classifier 3, Iteration: 0
	assign leaf[47] = !f[350] && !f[378] && !f[322] && !f[428];
	assign leaf[48] = !f[350] && !f[378] && !f[322] && f[428];
	assign leaf[49] = !f[350] && !f[378] && f[322] && !f[151];
	assign leaf[50] = !f[350] && !f[378] && f[322] && f[151];
	assign leaf[51] = !f[350] && f[378] && !f[176] && !f[592];
	assign leaf[52] = !f[350] && f[378] && !f[176] && f[592];
	assign leaf[53] = !f[350] && f[378] && f[176] && !f[543];
	assign leaf[54] = !f[350] && f[378] && f[176] && f[543];
	assign leaf[55] = f[350] && !f[489] && !f[290] && !f[179];
	assign leaf[56] = f[350] && !f[489] && !f[290] && f[179];
	assign leaf[57] = f[350] && !f[489] && f[290] && !f[318];
	assign leaf[58] = f[350] && !f[489] && f[290] && f[318];
	assign leaf[59] = f[350] && f[489] && !f[517] && !f[515];
	assign leaf[60] = f[350] && f[489] && !f[517] && f[515];
	assign leaf[61] = f[350] && f[489] && f[517] && !f[536];
	assign leaf[62] = f[350] && f[489] && f[517] && f[536];
	
	// Tree 4, Classifier 4, Iteration: 0
	assign leaf[63] = !f[211] && !f[428] && !f[402] && !f[398];
	assign leaf[64] = !f[211] && !f[428] && !f[402] && f[398];
	assign leaf[65] = !f[211] && !f[428] && f[402] && !f[155];
	assign leaf[66] = !f[211] && !f[428] && f[402] && f[155];
	assign leaf[67] = !f[211] && f[428] && !f[570] && !f[267];
	assign leaf[68] = !f[211] && f[428] && !f[570] && f[267];
	assign leaf[69] = !f[211] && f[428] && f[570] && !f[191];
	assign leaf[70] = !f[211] && f[428] && f[570] && f[191];
	assign leaf[71] = f[211] && !f[429] && !f[373] && !f[375];
	assign leaf[72] = f[211] && !f[429] && !f[373] && f[375];
	assign leaf[73] = f[211] && !f[429] && f[373] && !f[208];
	assign leaf[74] = f[211] && !f[429] && f[373] && f[208];
	assign leaf[75] = f[211] && f[429] && !f[210] && !f[600];
	assign leaf[76] = f[211] && f[429] && !f[210] && f[600];
	assign leaf[77] = f[211] && f[429] && f[210] && !f[213];
	assign leaf[78] = f[211] && f[429] && f[210] && f[213];
	
	// Tree 5, Classifier 5, Iteration: 0
	assign leaf[79] = !f[220] && !f[163] && !f[276] && !f[347];
	assign leaf[80] = !f[220] && !f[163] && !f[276] && f[347];
	assign leaf[81] = !f[220] && !f[163] && f[276] && !f[330];
	assign leaf[82] = !f[220] && !f[163] && f[276] && f[330];
	assign leaf[83] = !f[220] && f[163] && !f[272] && !f[302];
	assign leaf[84] = !f[220] && f[163] && !f[272] && f[302];
	assign leaf[85] = !f[220] && f[163] && f[272] && !f[299];
	assign leaf[86] = !f[220] && f[163] && f[272] && f[299];
	assign leaf[87] = f[220] && !f[328] && !f[358] && !f[326];
	assign leaf[88] = f[220] && !f[328] && !f[358] && f[326];
	assign leaf[89] = f[220] && !f[328] && f[358];
	assign leaf[90] = f[220] && f[328] && !f[355] && !f[276];
	assign leaf[91] = f[220] && f[328] && !f[355] && f[276];
	assign leaf[92] = f[220] && f[328] && f[355] && !f[382];
	assign leaf[93] = f[220] && f[328] && f[355] && f[382];
	
	// Tree 6, Classifier 6, Iteration: 0
	assign leaf[94] = !f[101] && !f[98] && !f[103] && !f[95];
	assign leaf[95] = !f[101] && !f[98] && !f[103] && f[95];
	assign leaf[96] = !f[101] && !f[98] && f[103] && !f[244];
	assign leaf[97] = !f[101] && !f[98] && f[103] && f[244];
	assign leaf[98] = !f[101] && f[98] && !f[213] && !f[267];
	assign leaf[99] = !f[101] && f[98] && !f[213] && f[267];
	assign leaf[100] = !f[101] && f[98] && f[213] && !f[291];
	assign leaf[101] = !f[101] && f[98] && f[213] && f[291];
	assign leaf[102] = f[101] && !f[243] && !f[594] && !f[269];
	assign leaf[103] = f[101] && !f[243] && !f[594] && f[269];
	assign leaf[104] = f[101] && !f[243] && f[594] && !f[292];
	assign leaf[105] = f[101] && !f[243] && f[594] && f[292];
	assign leaf[106] = f[101] && f[243] && !f[317] && !f[318];
	assign leaf[107] = f[101] && f[243] && !f[317] && f[318];
	assign leaf[108] = f[101] && f[243] && f[317] && !f[461];
	assign leaf[109] = f[101] && f[243] && f[317] && f[461];
	
	// Tree 7, Classifier 7, Iteration: 0
	assign leaf[110] = !f[739] && !f[742] && !f[709] && !f[712];
	assign leaf[111] = !f[739] && !f[742] && !f[709] && f[712];
	assign leaf[112] = !f[739] && !f[742] && f[709] && !f[405];
	assign leaf[113] = !f[739] && !f[742] && f[709] && f[405];
	assign leaf[114] = !f[739] && f[742] && !f[431] && !f[404];
	assign leaf[115] = !f[739] && f[742] && !f[431] && f[404];
	assign leaf[116] = !f[739] && f[742] && f[431] && !f[231];
	assign leaf[117] = !f[739] && f[742] && f[431] && f[231];
	assign leaf[118] = f[739] && !f[405] && !f[460] && !f[377];
	assign leaf[119] = f[739] && !f[405] && !f[460] && f[377];
	assign leaf[120] = f[739] && !f[405] && f[460] && !f[232];
	assign leaf[121] = f[739] && !f[405] && f[460] && f[232];
	assign leaf[122] = f[739] && f[405] && !f[233] && !f[207];
	assign leaf[123] = f[739] && f[405] && !f[233] && f[207];
	assign leaf[124] = f[739] && f[405] && f[233] && !f[374];
	assign leaf[125] = f[739] && f[405] && f[233] && f[374];
	
	// Tree 8, Classifier 8, Iteration: 0
	assign leaf[126] = !f[487] && !f[488] && !f[486] && !f[489];
	assign leaf[127] = !f[487] && !f[488] && !f[486] && f[489];
	assign leaf[128] = !f[487] && !f[488] && f[486] && !f[377];
	assign leaf[129] = !f[487] && !f[488] && f[486] && f[377];
	assign leaf[130] = !f[487] && f[488] && !f[659] && !f[376];
	assign leaf[131] = !f[487] && f[488] && !f[659] && f[376];
	assign leaf[132] = !f[487] && f[488] && f[659] && !f[347];
	assign leaf[133] = !f[487] && f[488] && f[659] && f[347];
	assign leaf[134] = f[487] && !f[656] && !f[276] && !f[657];
	assign leaf[135] = f[487] && !f[656] && !f[276] && f[657];
	assign leaf[136] = f[487] && !f[656] && f[276] && !f[214];
	assign leaf[137] = f[487] && !f[656] && f[276] && f[214];
	assign leaf[138] = f[487] && f[656] && !f[405] && !f[457];
	assign leaf[139] = f[487] && f[656] && !f[405] && f[457];
	assign leaf[140] = f[487] && f[656] && f[405] && !f[514];
	assign leaf[141] = f[487] && f[656] && f[405] && f[514];
	
	// Tree 9, Classifier 9, Iteration: 0
	assign leaf[142] = !f[717] && !f[713] && !f[715] && !f[711];
	assign leaf[143] = !f[717] && !f[713] && !f[715] && f[711];
	assign leaf[144] = !f[717] && !f[713] && f[715] && !f[210];
	assign leaf[145] = !f[717] && !f[713] && f[715] && f[210];
	assign leaf[146] = !f[717] && f[713] && !f[430] && !f[375];
	assign leaf[147] = !f[717] && f[713] && !f[430] && f[375];
	assign leaf[148] = !f[717] && f[713] && f[430] && !f[211];
	assign leaf[149] = !f[717] && f[713] && f[430] && f[211];
	assign leaf[150] = f[717] && !f[210] && !f[208] && !f[459];
	assign leaf[151] = f[717] && !f[210] && !f[208] && f[459];
	assign leaf[152] = f[717] && !f[210] && f[208] && !f[378];
	assign leaf[153] = f[717] && !f[210] && f[208] && f[378];
	assign leaf[154] = f[717] && f[210] && !f[231] && !f[685];
	assign leaf[155] = f[717] && f[210] && !f[231] && f[685];
	assign leaf[156] = f[717] && f[210] && f[231] && !f[398];
	assign leaf[157] = f[717] && f[210] && f[231] && f[398];
	
	// Tree 10, Classifier 0, Iteration: 1
	assign leaf[158] = !f[407] && !f[463] && !f[351] && !f[627];
	assign leaf[159] = !f[407] && !f[463] && !f[351] && f[627];
	assign leaf[160] = !f[407] && !f[463] && f[351] && !f[455];
	assign leaf[161] = !f[407] && !f[463] && f[351] && f[455];
	assign leaf[162] = !f[407] && f[463] && !f[321] && !f[415];
	assign leaf[163] = !f[407] && f[463] && !f[321] && f[415];
	assign leaf[164] = !f[407] && f[463] && f[321] && !f[511];
	assign leaf[165] = !f[407] && f[463] && f[321] && f[511];
	assign leaf[166] = f[407] && !f[359] && !f[512];
	assign leaf[167] = f[407] && !f[359] && f[512] && !f[322];
	assign leaf[168] = f[407] && !f[359] && f[512] && f[322];
	assign leaf[169] = f[407] && f[359] && !f[509] && !f[188];
	assign leaf[170] = f[407] && f[359] && !f[509] && f[188];
	assign leaf[171] = f[407] && f[359] && f[509] && !f[296];
	assign leaf[172] = f[407] && f[359] && f[509] && f[296];
	
	// Tree 11, Classifier 1, Iteration: 1
	assign leaf[173] = !f[409] && !f[378] && !f[379] && !f[377];
	assign leaf[174] = !f[409] && !f[378] && !f[379] && f[377];
	assign leaf[175] = !f[409] && !f[378] && f[379] && !f[353];
	assign leaf[176] = !f[409] && !f[378] && f[379] && f[353];
	assign leaf[177] = !f[409] && f[378] && !f[550] && !f[319];
	assign leaf[178] = !f[409] && f[378] && !f[550] && f[319];
	assign leaf[179] = !f[409] && f[378] && f[550] && !f[293];
	assign leaf[180] = !f[409] && f[378] && f[550] && f[293];
	assign leaf[181] = f[409] && !f[410] && !f[323] && !f[594];
	assign leaf[182] = f[409] && !f[410] && !f[323] && f[594];
	assign leaf[183] = f[409] && !f[410] && f[323] && !f[544];
	assign leaf[184] = f[409] && !f[410] && f[323] && f[544];
	assign leaf[185] = f[409] && f[410] && !f[171] && !f[613];
	assign leaf[186] = f[409] && f[410] && !f[171] && f[613];
	assign leaf[187] = f[409] && f[410] && f[171];
	
	// Tree 12, Classifier 2, Iteration: 1
	assign leaf[188] = !f[542] && !f[512] && !f[99] && !f[571];
	assign leaf[189] = !f[542] && !f[512] && !f[99] && f[571];
	assign leaf[190] = !f[542] && !f[512] && f[99] && !f[482];
	assign leaf[191] = !f[542] && !f[512] && f[99] && f[482];
	assign leaf[192] = !f[542] && f[512] && !f[346] && !f[658];
	assign leaf[193] = !f[542] && f[512] && !f[346] && f[658];
	assign leaf[194] = !f[542] && f[512] && f[346] && !f[97];
	assign leaf[195] = !f[542] && f[512] && f[346] && f[97];
	assign leaf[196] = f[542] && !f[347] && !f[344] && !f[350];
	assign leaf[197] = f[542] && !f[347] && !f[344] && f[350];
	assign leaf[198] = f[542] && !f[347] && f[344] && !f[372];
	assign leaf[199] = f[542] && !f[347] && f[344] && f[372];
	assign leaf[200] = f[542] && f[347] && !f[528] && !f[582];
	assign leaf[201] = f[542] && f[347] && !f[528] && f[582];
	assign leaf[202] = f[542] && f[347] && f[528] && !f[414];
	assign leaf[203] = f[542] && f[347] && f[528] && f[414];
	
	// Tree 13, Classifier 3, Iteration: 1
	assign leaf[204] = !f[151] && !f[622] && !f[179] && !f[564];
	assign leaf[205] = !f[151] && !f[622] && !f[179] && f[564];
	assign leaf[206] = !f[151] && !f[622] && f[179] && !f[317];
	assign leaf[207] = !f[151] && !f[622] && f[179] && f[317];
	assign leaf[208] = !f[151] && f[622] && !f[351] && !f[379];
	assign leaf[209] = !f[151] && f[622] && !f[351] && f[379];
	assign leaf[210] = !f[151] && f[622] && f[351] && !f[486];
	assign leaf[211] = !f[151] && f[622] && f[351] && f[486];
	assign leaf[212] = f[151] && !f[514] && !f[289] && !f[518];
	assign leaf[213] = f[151] && !f[514] && !f[289] && f[518];
	assign leaf[214] = f[151] && !f[514] && f[289] && !f[267];
	assign leaf[215] = f[151] && !f[514] && f[289] && f[267];
	assign leaf[216] = f[151] && f[514] && !f[321] && !f[679];
	assign leaf[217] = f[151] && f[514] && !f[321] && f[679];
	assign leaf[218] = f[151] && f[514] && f[321] && !f[459];
	assign leaf[219] = f[151] && f[514] && f[321] && f[459];
	
	// Tree 14, Classifier 4, Iteration: 1
	assign leaf[220] = !f[400] && !f[402] && !f[398] && !f[375];
	assign leaf[221] = !f[400] && !f[402] && !f[398] && f[375];
	assign leaf[222] = !f[400] && !f[402] && f[398] && !f[458];
	assign leaf[223] = !f[400] && !f[402] && f[398] && f[458];
	assign leaf[224] = !f[400] && f[402] && !f[183] && !f[239];
	assign leaf[225] = !f[400] && f[402] && !f[183] && f[239];
	assign leaf[226] = !f[400] && f[402] && f[183] && !f[185];
	assign leaf[227] = !f[400] && f[402] && f[183] && f[185];
	assign leaf[228] = f[400] && !f[210] && !f[154] && !f[266];
	assign leaf[229] = f[400] && !f[210] && !f[154] && f[266];
	assign leaf[230] = f[400] && !f[210] && f[154] && !f[155];
	assign leaf[231] = f[400] && !f[210] && f[154] && f[155];
	assign leaf[232] = f[400] && f[210] && !f[463] && !f[628];
	assign leaf[233] = f[400] && f[210] && !f[463] && f[628];
	assign leaf[234] = f[400] && f[210] && f[463] && !f[212];
	assign leaf[235] = f[400] && f[210] && f[463] && f[212];
	
	// Tree 15, Classifier 5, Iteration: 1
	assign leaf[236] = !f[347] && !f[248] && !f[192] && !f[375];
	assign leaf[237] = !f[347] && !f[248] && !f[192] && f[375];
	assign leaf[238] = !f[347] && !f[248] && f[192] && !f[300];
	assign leaf[239] = !f[347] && !f[248] && f[192] && f[300];
	assign leaf[240] = !f[347] && f[248] && !f[355] && !f[359];
	assign leaf[241] = !f[347] && f[248] && !f[355] && f[359];
	assign leaf[242] = !f[347] && f[248] && f[355];
	assign leaf[243] = f[347] && !f[326] && !f[515] && !f[329];
	assign leaf[244] = f[347] && !f[326] && !f[515] && f[329];
	assign leaf[245] = f[347] && !f[326] && f[515] && !f[247];
	assign leaf[246] = f[347] && !f[326] && f[515] && f[247];
	assign leaf[247] = f[347] && f[326] && !f[408] && !f[270];
	assign leaf[248] = f[347] && f[326] && !f[408] && f[270];
	assign leaf[249] = f[347] && f[326] && f[408] && !f[304];
	assign leaf[250] = f[347] && f[326] && f[408] && f[304];
	
	// Tree 16, Classifier 6, Iteration: 1
	assign leaf[251] = !f[514] && !f[101] && !f[70] && !f[105];
	assign leaf[252] = !f[514] && !f[101] && !f[70] && f[105];
	assign leaf[253] = !f[514] && !f[101] && f[70] && !f[156];
	assign leaf[254] = !f[514] && !f[101] && f[70] && f[156];
	assign leaf[255] = !f[514] && f[101] && !f[625] && !f[237];
	assign leaf[256] = !f[514] && f[101] && !f[625] && f[237];
	assign leaf[257] = !f[514] && f[101] && f[625] && !f[414];
	assign leaf[258] = !f[514] && f[101] && f[625] && f[414];
	assign leaf[259] = f[514] && !f[242] && !f[245] && !f[268];
	assign leaf[260] = f[514] && !f[242] && !f[245] && f[268];
	assign leaf[261] = f[514] && !f[242] && f[245] && !f[120];
	assign leaf[262] = f[514] && !f[242] && f[245] && f[120];
	assign leaf[263] = f[514] && f[242] && !f[105] && !f[135];
	assign leaf[264] = f[514] && f[242] && !f[105] && f[135];
	assign leaf[265] = f[514] && f[242] && f[105] && !f[325];
	assign leaf[266] = f[514] && f[242] && f[105] && f[325];
	
	// Tree 17, Classifier 7, Iteration: 1
	assign leaf[267] = !f[405] && !f[155] && !f[457] && !f[568];
	assign leaf[268] = !f[405] && !f[155] && !f[457] && f[568];
	assign leaf[269] = !f[405] && !f[155] && f[457] && !f[229];
	assign leaf[270] = !f[405] && !f[155] && f[457] && f[229];
	assign leaf[271] = !f[405] && f[155] && !f[678] && !f[578];
	assign leaf[272] = !f[405] && f[155] && !f[678] && f[578];
	assign leaf[273] = !f[405] && f[155] && f[678] && !f[603];
	assign leaf[274] = !f[405] && f[155] && f[678] && f[603];
	assign leaf[275] = f[405] && !f[231] && !f[708] && !f[710];
	assign leaf[276] = f[405] && !f[231] && !f[708] && f[710];
	assign leaf[277] = f[405] && !f[231] && f[708] && !f[542];
	assign leaf[278] = f[405] && !f[231] && f[708] && f[542];
	assign leaf[279] = f[405] && f[231] && !f[606] && !f[264];
	assign leaf[280] = f[405] && f[231] && !f[606] && f[264];
	assign leaf[281] = f[405] && f[231] && f[606] && !f[312];
	assign leaf[282] = f[405] && f[231] && f[606] && f[312];
	
	// Tree 18, Classifier 8, Iteration: 1
	assign leaf[283] = !f[376] && !f[349] && !f[403] && !f[276];
	assign leaf[284] = !f[376] && !f[349] && !f[403] && f[276];
	assign leaf[285] = !f[376] && !f[349] && f[403] && !f[515];
	assign leaf[286] = !f[376] && !f[349] && f[403] && f[515];
	assign leaf[287] = !f[376] && f[349] && !f[295] && !f[460];
	assign leaf[288] = !f[376] && f[349] && !f[295] && f[460];
	assign leaf[289] = !f[376] && f[349] && f[295] && !f[459];
	assign leaf[290] = !f[376] && f[349] && f[295] && f[459];
	assign leaf[291] = f[376] && !f[461] && !f[486] && !f[485];
	assign leaf[292] = f[376] && !f[461] && !f[486] && f[485];
	assign leaf[293] = f[376] && !f[461] && f[486] && !f[407];
	assign leaf[294] = f[376] && !f[461] && f[486] && f[407];
	assign leaf[295] = f[376] && f[461] && !f[657] && !f[623];
	assign leaf[296] = f[376] && f[461] && !f[657] && f[623];
	assign leaf[297] = f[376] && f[461] && f[657] && !f[515];
	assign leaf[298] = f[376] && f[461] && f[657] && f[515];
	
	// Tree 19, Classifier 9, Iteration: 1
	assign leaf[299] = !f[156] && !f[211] && !f[720] && !f[239];
	assign leaf[300] = !f[156] && !f[211] && !f[720] && f[239];
	assign leaf[301] = !f[156] && !f[211] && f[720] && !f[209];
	assign leaf[302] = !f[156] && !f[211] && f[720] && f[209];
	assign leaf[303] = !f[156] && f[211] && !f[409] && !f[408];
	assign leaf[304] = !f[156] && f[211] && !f[409] && f[408];
	assign leaf[305] = !f[156] && f[211] && f[409] && !f[345];
	assign leaf[306] = !f[156] && f[211] && f[409] && f[345];
	assign leaf[307] = f[156] && !f[128] && !f[409] && !f[439];
	assign leaf[308] = f[156] && !f[128] && !f[409] && f[439];
	assign leaf[309] = f[156] && !f[128] && f[409] && !f[626];
	assign leaf[310] = f[156] && !f[128] && f[409] && f[626];
	assign leaf[311] = f[156] && f[128] && !f[368];
	assign leaf[312] = f[156] && f[128] && f[368];
	
	// Tree 20, Classifier 0, Iteration: 2
	assign leaf[313] = !f[407] && !f[490] && !f[352] && !f[184];
	assign leaf[314] = !f[407] && !f[490] && !f[352] && f[184];
	assign leaf[315] = !f[407] && !f[490] && f[352] && !f[456];
	assign leaf[316] = !f[407] && !f[490] && f[352] && f[456];
	assign leaf[317] = !f[407] && f[490] && !f[359] && !f[347];
	assign leaf[318] = !f[407] && f[490] && !f[359] && f[347];
	assign leaf[319] = !f[407] && f[490] && f[359] && !f[453];
	assign leaf[320] = !f[407] && f[490] && f[359] && f[453];
	assign leaf[321] = f[407] && !f[359] && !f[512];
	assign leaf[322] = f[407] && !f[359] && f[512] && !f[294];
	assign leaf[323] = f[407] && !f[359] && f[512] && f[294];
	assign leaf[324] = f[407] && f[359] && !f[322] && !f[187];
	assign leaf[325] = f[407] && f[359] && !f[322] && f[187];
	assign leaf[326] = f[407] && f[359] && f[322] && !f[432];
	assign leaf[327] = f[407] && f[359] && f[322] && f[432];
	
	// Tree 21, Classifier 1, Iteration: 2
	assign leaf[328] = !f[437] && !f[262] && !f[406] && !f[407];
	assign leaf[329] = !f[437] && !f[262] && !f[406] && f[407];
	assign leaf[330] = !f[437] && !f[262] && f[406] && !f[178];
	assign leaf[331] = !f[437] && !f[262] && f[406] && f[178];
	assign leaf[332] = !f[437] && f[262] && !f[325] && !f[350];
	assign leaf[333] = !f[437] && f[262] && !f[325] && f[350];
	assign leaf[334] = !f[437] && f[262] && f[325];
	assign leaf[335] = f[437] && !f[438] && !f[322] && !f[622];
	assign leaf[336] = f[437] && !f[438] && !f[322] && f[622];
	assign leaf[337] = f[437] && !f[438] && f[322] && !f[545];
	assign leaf[338] = f[437] && !f[438] && f[322] && f[545];
	assign leaf[339] = f[437] && f[438] && !f[613] && !f[69];
	assign leaf[340] = f[437] && f[438] && !f[613] && f[69];
	assign leaf[341] = f[437] && f[438] && f[613];
	
	// Tree 22, Classifier 2, Iteration: 2
	assign leaf[342] = !f[568] && !f[123] && !f[539] && !f[473];
	assign leaf[343] = !f[568] && !f[123] && !f[539] && f[473];
	assign leaf[344] = !f[568] && !f[123] && f[539] && !f[346];
	assign leaf[345] = !f[568] && !f[123] && f[539] && f[346];
	assign leaf[346] = !f[568] && f[123] && !f[345] && !f[348];
	assign leaf[347] = !f[568] && f[123] && !f[345] && f[348];
	assign leaf[348] = !f[568] && f[123] && f[345] && !f[664];
	assign leaf[349] = !f[568] && f[123] && f[345] && f[664];
	assign leaf[350] = f[568] && !f[517] && !f[460] && !f[98];
	assign leaf[351] = f[568] && !f[517] && !f[460] && f[98];
	assign leaf[352] = f[568] && !f[517] && f[460] && !f[348];
	assign leaf[353] = f[568] && !f[517] && f[460] && f[348];
	assign leaf[354] = f[568] && f[517] && !f[320] && !f[156];
	assign leaf[355] = f[568] && f[517] && !f[320] && f[156];
	assign leaf[356] = f[568] && f[517] && f[320] && !f[580];
	assign leaf[357] = f[568] && f[517] && f[320] && f[580];
	
	// Tree 23, Classifier 3, Iteration: 2
	assign leaf[358] = !f[350] && !f[378] && !f[322] && !f[406];
	assign leaf[359] = !f[350] && !f[378] && !f[322] && f[406];
	assign leaf[360] = !f[350] && !f[378] && f[322] && !f[153];
	assign leaf[361] = !f[350] && !f[378] && f[322] && f[153];
	assign leaf[362] = !f[350] && f[378] && !f[318] && !f[543];
	assign leaf[363] = !f[350] && f[378] && !f[318] && f[543];
	assign leaf[364] = !f[350] && f[378] && f[318] && !f[148];
	assign leaf[365] = !f[350] && f[378] && f[318] && f[148];
	assign leaf[366] = f[350] && !f[517] && !f[487] && !f[316];
	assign leaf[367] = f[350] && !f[517] && !f[487] && f[316];
	assign leaf[368] = f[350] && !f[517] && f[487] && !f[542];
	assign leaf[369] = f[350] && !f[517] && f[487] && f[542];
	assign leaf[370] = f[350] && f[517] && !f[462] && !f[410];
	assign leaf[371] = f[350] && f[517] && !f[462] && f[410];
	assign leaf[372] = f[350] && f[517] && f[462] && !f[594];
	assign leaf[373] = f[350] && f[517] && f[462] && f[594];
	
	// Tree 24, Classifier 4, Iteration: 2
	assign leaf[374] = !f[183] && !f[267] && !f[437] && !f[464];
	assign leaf[375] = !f[183] && !f[267] && !f[437] && f[464];
	assign leaf[376] = !f[183] && !f[267] && f[437] && !f[126];
	assign leaf[377] = !f[183] && !f[267] && f[437] && f[126];
	assign leaf[378] = !f[183] && f[267] && !f[429] && !f[375];
	assign leaf[379] = !f[183] && f[267] && !f[429] && f[375];
	assign leaf[380] = !f[183] && f[267] && f[429] && !f[237];
	assign leaf[381] = !f[183] && f[267] && f[429] && f[237];
	assign leaf[382] = f[183] && !f[180] && !f[662] && !f[464];
	assign leaf[383] = f[183] && !f[180] && !f[662] && f[464];
	assign leaf[384] = f[183] && !f[180] && f[662] && !f[235];
	assign leaf[385] = f[183] && !f[180] && f[662] && f[235];
	assign leaf[386] = f[183] && f[180] && !f[182] && !f[153];
	assign leaf[387] = f[183] && f[180] && !f[182] && f[153];
	assign leaf[388] = f[183] && f[180] && f[182] && !f[184];
	assign leaf[389] = f[183] && f[180] && f[182] && f[184];
	
	// Tree 25, Classifier 5, Iteration: 2
	assign leaf[390] = !f[326] && !f[296] && !f[356] && !f[655];
	assign leaf[391] = !f[326] && !f[296] && !f[356] && f[655];
	assign leaf[392] = !f[326] && !f[296] && f[356] && !f[351];
	assign leaf[393] = !f[326] && !f[296] && f[356] && f[351];
	assign leaf[394] = !f[326] && f[296] && !f[246] && !f[275];
	assign leaf[395] = !f[326] && f[296] && !f[246] && f[275];
	assign leaf[396] = !f[326] && f[296] && f[246] && !f[357];
	assign leaf[397] = !f[326] && f[296] && f[246] && f[357];
	assign leaf[398] = f[326] && !f[304] && !f[322] && !f[332];
	assign leaf[399] = f[326] && !f[304] && !f[322] && f[332];
	assign leaf[400] = f[326] && !f[304] && f[322] && !f[298];
	assign leaf[401] = f[326] && !f[304] && f[322] && f[298];
	assign leaf[402] = f[326] && f[304] && !f[381] && !f[215];
	assign leaf[403] = f[326] && f[304] && !f[381] && f[215];
	assign leaf[404] = f[326] && f[304] && f[381] && !f[322];
	assign leaf[405] = f[326] && f[304] && f[381] && f[322];
	
	// Tree 26, Classifier 6, Iteration: 2
	assign leaf[406] = !f[543] && !f[104] && !f[101] && !f[69];
	assign leaf[407] = !f[543] && !f[104] && !f[101] && f[69];
	assign leaf[408] = !f[543] && !f[104] && f[101] && !f[402];
	assign leaf[409] = !f[543] && !f[104] && f[101] && f[402];
	assign leaf[410] = !f[543] && f[104] && !f[541] && !f[266];
	assign leaf[411] = !f[543] && f[104] && !f[541] && f[266];
	assign leaf[412] = !f[543] && f[104] && f[541] && !f[103];
	assign leaf[413] = !f[543] && f[104] && f[541] && f[103];
	assign leaf[414] = f[543] && !f[242] && !f[655] && !f[216];
	assign leaf[415] = f[543] && !f[242] && !f[655] && f[216];
	assign leaf[416] = f[543] && !f[242] && f[655] && !f[131];
	assign leaf[417] = f[543] && !f[242] && f[655] && f[131];
	assign leaf[418] = f[543] && f[242] && !f[106] && !f[104];
	assign leaf[419] = f[543] && f[242] && !f[106] && f[104];
	assign leaf[420] = f[543] && f[242] && f[106] && !f[325];
	assign leaf[421] = f[543] && f[242] && f[106] && f[325];
	
	// Tree 27, Classifier 7, Iteration: 2
	assign leaf[422] = !f[405] && !f[156] && !f[458] && !f[153];
	assign leaf[423] = !f[405] && !f[156] && !f[458] && f[153];
	assign leaf[424] = !f[405] && !f[156] && f[458] && !f[231];
	assign leaf[425] = !f[405] && !f[156] && f[458] && f[231];
	assign leaf[426] = !f[405] && f[156] && !f[678] && !f[597];
	assign leaf[427] = !f[405] && f[156] && !f[678] && f[597];
	assign leaf[428] = !f[405] && f[156] && f[678] && !f[570];
	assign leaf[429] = !f[405] && f[156] && f[678] && f[570];
	assign leaf[430] = f[405] && !f[231] && !f[257] && !f[705];
	assign leaf[431] = f[405] && !f[231] && !f[257] && f[705];
	assign leaf[432] = f[405] && !f[231] && f[257] && !f[289];
	assign leaf[433] = f[405] && !f[231] && f[257] && f[289];
	assign leaf[434] = f[405] && f[231] && !f[519] && !f[500];
	assign leaf[435] = f[405] && f[231] && !f[519] && f[500];
	assign leaf[436] = f[405] && f[231] && f[519] && !f[550];
	assign leaf[437] = f[405] && f[231] && f[519] && f[550];
	
	// Tree 28, Classifier 8, Iteration: 2
	assign leaf[438] = !f[657] && !f[275] && !f[376] && !f[629];
	assign leaf[439] = !f[657] && !f[275] && !f[376] && f[629];
	assign leaf[440] = !f[657] && !f[275] && f[376] && !f[662];
	assign leaf[441] = !f[657] && !f[275] && f[376] && f[662];
	assign leaf[442] = !f[657] && f[275] && !f[486] && !f[488];
	assign leaf[443] = !f[657] && f[275] && !f[486] && f[488];
	assign leaf[444] = !f[657] && f[275] && f[486] && !f[466];
	assign leaf[445] = !f[657] && f[275] && f[486] && f[466];
	assign leaf[446] = f[657] && !f[515] && !f[513] && !f[516];
	assign leaf[447] = f[657] && !f[515] && !f[513] && f[516];
	assign leaf[448] = f[657] && !f[515] && f[513] && !f[404];
	assign leaf[449] = f[657] && !f[515] && f[513] && f[404];
	assign leaf[450] = f[657] && f[515] && !f[433] && !f[378];
	assign leaf[451] = f[657] && f[515] && !f[433] && f[378];
	assign leaf[452] = f[657] && f[515] && f[433] && !f[573];
	assign leaf[453] = f[657] && f[515] && f[433] && f[573];
	
	// Tree 29, Classifier 9, Iteration: 2
	assign leaf[454] = !f[597] && !f[381] && !f[721] && !f[383];
	assign leaf[455] = !f[597] && !f[381] && !f[721] && f[383];
	assign leaf[456] = !f[597] && !f[381] && f[721] && !f[488];
	assign leaf[457] = !f[597] && !f[381] && f[721] && f[488];
	assign leaf[458] = !f[597] && f[381] && !f[211] && !f[238];
	assign leaf[459] = !f[597] && f[381] && !f[211] && f[238];
	assign leaf[460] = !f[597] && f[381] && f[211] && !f[205];
	assign leaf[461] = !f[597] && f[381] && f[211] && f[205];
	assign leaf[462] = f[597] && !f[707] && !f[706] && !f[708];
	assign leaf[463] = f[597] && !f[707] && !f[706] && f[708];
	assign leaf[464] = f[597] && !f[707] && f[706];
	assign leaf[465] = f[597] && f[707] && !f[376] && !f[429];
	assign leaf[466] = f[597] && f[707] && !f[376] && f[429];
	assign leaf[467] = f[597] && f[707] && f[376] && !f[219];
	assign leaf[468] = f[597] && f[707] && f[376] && f[219];
	
	// Tree 30, Classifier 0, Iteration: 3
	assign leaf[469] = !f[434] && !f[380] && !f[489] && !f[484];
	assign leaf[470] = !f[434] && !f[380] && !f[489] && f[484];
	assign leaf[471] = !f[434] && !f[380] && f[489] && !f[386];
	assign leaf[472] = !f[434] && !f[380] && f[489] && f[386];
	assign leaf[473] = !f[434] && f[380] && !f[513] && !f[331];
	assign leaf[474] = !f[434] && f[380] && !f[513] && f[331];
	assign leaf[475] = !f[434] && f[380] && f[513] && !f[267];
	assign leaf[476] = !f[434] && f[380] && f[513] && f[267];
	assign leaf[477] = f[434] && !f[386] && !f[387];
	assign leaf[478] = f[434] && !f[386] && f[387] && !f[209];
	assign leaf[479] = f[434] && !f[386] && f[387] && f[209];
	assign leaf[480] = f[434] && f[386] && !f[625] && !f[219];
	assign leaf[481] = f[434] && f[386] && !f[625] && f[219];
	assign leaf[482] = f[434] && f[386] && f[625] && !f[468];
	assign leaf[483] = f[434] && f[386] && f[625] && f[468];
	
	// Tree 31, Classifier 1, Iteration: 3
	assign leaf[484] = !f[350] && !f[351] && !f[382] && !f[374];
	assign leaf[485] = !f[350] && !f[351] && !f[382] && f[374];
	assign leaf[486] = !f[350] && !f[351] && f[382];
	assign leaf[487] = !f[350] && f[351] && !f[209] && !f[431];
	assign leaf[488] = !f[350] && f[351] && !f[209] && f[431];
	assign leaf[489] = !f[350] && f[351] && f[209] && !f[406];
	assign leaf[490] = !f[350] && f[351] && f[209] && f[406];
	assign leaf[491] = f[350] && !f[375] && !f[234] && !f[327];
	assign leaf[492] = f[350] && !f[375] && !f[234] && f[327];
	assign leaf[493] = f[350] && !f[375] && f[234] && !f[297];
	assign leaf[494] = f[350] && !f[375] && f[234] && f[297];
	assign leaf[495] = f[350] && f[375] && !f[374] && !f[517];
	assign leaf[496] = f[350] && f[375] && !f[374] && f[517];
	assign leaf[497] = f[350] && f[375] && f[374] && !f[294];
	assign leaf[498] = f[350] && f[375] && f[374] && f[294];
	
	// Tree 32, Classifier 2, Iteration: 3
	assign leaf[499] = !f[346] && !f[569] && !f[511] && !f[582];
	assign leaf[500] = !f[346] && !f[569] && !f[511] && f[582];
	assign leaf[501] = !f[346] && !f[569] && f[511] && !f[343];
	assign leaf[502] = !f[346] && !f[569] && f[511] && f[343];
	assign leaf[503] = !f[346] && f[569] && !f[321] && !f[371];
	assign leaf[504] = !f[346] && f[569] && !f[321] && f[371];
	assign leaf[505] = !f[346] && f[569] && f[321] && !f[554];
	assign leaf[506] = !f[346] && f[569] && f[321] && f[554];
	assign leaf[507] = f[346] && !f[528] && !f[584] && !f[637];
	assign leaf[508] = f[346] && !f[528] && !f[584] && f[637];
	assign leaf[509] = f[346] && !f[528] && f[584];
	assign leaf[510] = f[346] && f[528] && !f[413] && !f[551];
	assign leaf[511] = f[346] && f[528] && !f[413] && f[551];
	assign leaf[512] = f[346] && f[528] && f[413] && !f[493];
	assign leaf[513] = f[346] && f[528] && f[413] && f[493];
	
	// Tree 33, Classifier 3, Iteration: 3
	assign leaf[514] = !f[490] && !f[317] && !f[487] && !f[291];
	assign leaf[515] = !f[490] && !f[317] && !f[487] && f[291];
	assign leaf[516] = !f[490] && !f[317] && f[487] && !f[515];
	assign leaf[517] = !f[490] && !f[317] && f[487] && f[515];
	assign leaf[518] = !f[490] && f[317] && !f[147] && !f[322];
	assign leaf[519] = !f[490] && f[317] && !f[147] && f[322];
	assign leaf[520] = !f[490] && f[317] && f[147] && !f[259];
	assign leaf[521] = !f[490] && f[317] && f[147] && f[259];
	assign leaf[522] = f[490] && !f[178] && !f[649] && !f[297];
	assign leaf[523] = f[490] && !f[178] && !f[649] && f[297];
	assign leaf[524] = f[490] && !f[178] && f[649] && !f[515];
	assign leaf[525] = f[490] && !f[178] && f[649] && f[515];
	assign leaf[526] = f[490] && f[178] && !f[657] && !f[714];
	assign leaf[527] = f[490] && f[178] && !f[657] && f[714];
	assign leaf[528] = f[490] && f[178] && f[657] && !f[545];
	assign leaf[529] = f[490] && f[178] && f[657] && f[545];
	
	// Tree 34, Classifier 4, Iteration: 3
	assign leaf[530] = !f[401] && !f[399] && !f[374] && !f[397];
	assign leaf[531] = !f[401] && !f[399] && !f[374] && f[397];
	assign leaf[532] = !f[401] && !f[399] && f[374] && !f[184];
	assign leaf[533] = !f[401] && !f[399] && f[374] && f[184];
	assign leaf[534] = !f[401] && f[399] && !f[458] && !f[487];
	assign leaf[535] = !f[401] && f[399] && !f[458] && f[487];
	assign leaf[536] = !f[401] && f[399] && f[458] && !f[210];
	assign leaf[537] = !f[401] && f[399] && f[458] && f[210];
	assign leaf[538] = f[401] && !f[569] && !f[463] && !f[210];
	assign leaf[539] = f[401] && !f[569] && !f[463] && f[210];
	assign leaf[540] = f[401] && !f[569] && f[463] && !f[209];
	assign leaf[541] = f[401] && !f[569] && f[463] && f[209];
	assign leaf[542] = f[401] && f[569] && !f[488] && !f[136];
	assign leaf[543] = f[401] && f[569] && !f[488] && f[136];
	assign leaf[544] = f[401] && f[569] && f[488] && !f[574];
	assign leaf[545] = f[401] && f[569] && f[488] && f[574];
	
	// Tree 35, Classifier 5, Iteration: 3
	assign leaf[546] = !f[489] && !f[298] && !f[300] && !f[295];
	assign leaf[547] = !f[489] && !f[298] && !f[300] && f[295];
	assign leaf[548] = !f[489] && !f[298] && f[300] && !f[328];
	assign leaf[549] = !f[489] && !f[298] && f[300] && f[328];
	assign leaf[550] = !f[489] && f[298] && !f[275] && !f[219];
	assign leaf[551] = !f[489] && f[298] && !f[275] && f[219];
	assign leaf[552] = !f[489] && f[298] && f[275] && !f[357];
	assign leaf[553] = !f[489] && f[298] && f[275] && f[357];
	assign leaf[554] = f[489] && !f[248] && !f[407] && !f[437];
	assign leaf[555] = f[489] && !f[248] && !f[407] && f[437];
	assign leaf[556] = f[489] && !f[248] && f[407] && !f[276];
	assign leaf[557] = f[489] && !f[248] && f[407] && f[276];
	assign leaf[558] = f[489] && f[248] && !f[355] && !f[385];
	assign leaf[559] = f[489] && f[248] && !f[355] && f[385];
	assign leaf[560] = f[489] && f[248] && f[355] && !f[323];
	assign leaf[561] = f[489] && f[248] && f[355] && f[323];
	
	// Tree 36, Classifier 6, Iteration: 3
	assign leaf[562] = !f[543] && !f[570] && !f[68] && !f[70];
	assign leaf[563] = !f[543] && !f[570] && !f[68] && f[70];
	assign leaf[564] = !f[543] && !f[570] && f[68];
	assign leaf[565] = !f[543] && f[570] && !f[271] && !f[457];
	assign leaf[566] = !f[543] && f[570] && !f[271] && f[457];
	assign leaf[567] = !f[543] && f[570] && f[271] && !f[92];
	assign leaf[568] = !f[543] && f[570] && f[271] && f[92];
	assign leaf[569] = f[543] && !f[242] && !f[575] && !f[296];
	assign leaf[570] = f[543] && !f[242] && !f[575] && f[296];
	assign leaf[571] = f[543] && !f[242] && f[575] && !f[625];
	assign leaf[572] = f[543] && !f[242] && f[575] && f[625];
	assign leaf[573] = f[543] && f[242] && !f[105] && !f[457];
	assign leaf[574] = f[543] && f[242] && !f[105] && f[457];
	assign leaf[575] = f[543] && f[242] && f[105] && !f[298];
	assign leaf[576] = f[543] && f[242] && f[105] && f[298];
	
	// Tree 37, Classifier 7, Iteration: 3
	assign leaf[577] = !f[405] && !f[268] && !f[430] && !f[154];
	assign leaf[578] = !f[405] && !f[268] && !f[430] && f[154];
	assign leaf[579] = !f[405] && !f[268] && f[430] && !f[256];
	assign leaf[580] = !f[405] && !f[268] && f[430] && f[256];
	assign leaf[581] = !f[405] && f[268] && !f[156] && !f[430];
	assign leaf[582] = !f[405] && f[268] && !f[156] && f[430];
	assign leaf[583] = !f[405] && f[268] && f[156] && !f[490];
	assign leaf[584] = !f[405] && f[268] && f[156] && f[490];
	assign leaf[585] = f[405] && !f[268] && !f[707] && !f[312];
	assign leaf[586] = f[405] && !f[268] && !f[707] && f[312];
	assign leaf[587] = f[405] && !f[268] && f[707] && !f[515];
	assign leaf[588] = f[405] && !f[268] && f[707] && f[515];
	assign leaf[589] = f[405] && f[268] && !f[235] && !f[285];
	assign leaf[590] = f[405] && f[268] && !f[235] && f[285];
	assign leaf[591] = f[405] && f[268] && f[235] && !f[376];
	assign leaf[592] = f[405] && f[268] && f[235] && f[376];
	
	// Tree 38, Classifier 8, Iteration: 3
	assign leaf[593] = !f[405] && !f[432] && !f[378] && !f[460];
	assign leaf[594] = !f[405] && !f[432] && !f[378] && f[460];
	assign leaf[595] = !f[405] && !f[432] && f[378] && !f[488];
	assign leaf[596] = !f[405] && !f[432] && f[378] && f[488];
	assign leaf[597] = !f[405] && f[432] && !f[457] && !f[516];
	assign leaf[598] = !f[405] && f[432] && !f[457] && f[516];
	assign leaf[599] = !f[405] && f[432] && f[457] && !f[332];
	assign leaf[600] = !f[405] && f[432] && f[457] && f[332];
	assign leaf[601] = f[405] && !f[300] && !f[319] && !f[346];
	assign leaf[602] = f[405] && !f[300] && !f[319] && f[346];
	assign leaf[603] = f[405] && !f[300] && f[319] && !f[402];
	assign leaf[604] = f[405] && !f[300] && f[319] && f[402];
	assign leaf[605] = f[405] && f[300] && !f[438] && !f[183];
	assign leaf[606] = f[405] && f[300] && !f[438] && f[183];
	assign leaf[607] = f[405] && f[300] && f[438] && !f[660];
	assign leaf[608] = f[405] && f[300] && f[438] && f[660];
	
	// Tree 39, Classifier 9, Iteration: 3
	assign leaf[609] = !f[569] && !f[381] && !f[342] && !f[290];
	assign leaf[610] = !f[569] && !f[381] && !f[342] && f[290];
	assign leaf[611] = !f[569] && !f[381] && f[342] && !f[209];
	assign leaf[612] = !f[569] && !f[381] && f[342] && f[209];
	assign leaf[613] = !f[569] && f[381] && !f[211] && !f[239];
	assign leaf[614] = !f[569] && f[381] && !f[211] && f[239];
	assign leaf[615] = !f[569] && f[381] && f[211] && !f[155];
	assign leaf[616] = !f[569] && f[381] && f[211] && f[155];
	assign leaf[617] = f[569] && !f[692] && !f[706] && !f[707];
	assign leaf[618] = f[569] && !f[692] && !f[706] && f[707];
	assign leaf[619] = f[569] && !f[692] && f[706] && !f[377];
	assign leaf[620] = f[569] && !f[692] && f[706] && f[377];
	assign leaf[621] = f[569] && f[692] && !f[482] && !f[511];
	assign leaf[622] = f[569] && f[692] && !f[482] && f[511];
	assign leaf[623] = f[569] && f[692] && f[482];
	
	// Tree 40, Classifier 0, Iteration: 4
	assign leaf[624] = !f[407] && !f[511] && !f[513] && !f[481];
	assign leaf[625] = !f[407] && !f[511] && !f[513] && f[481];
	assign leaf[626] = !f[407] && !f[511] && f[513] && !f[490];
	assign leaf[627] = !f[407] && !f[511] && f[513] && f[490];
	assign leaf[628] = !f[407] && f[511] && !f[488] && !f[379];
	assign leaf[629] = !f[407] && f[511] && !f[488] && f[379];
	assign leaf[630] = !f[407] && f[511] && f[488] && !f[400];
	assign leaf[631] = !f[407] && f[511] && f[488] && f[400];
	assign leaf[632] = f[407] && !f[359] && !f[512] && !f[396];
	assign leaf[633] = f[407] && !f[359] && !f[512] && f[396];
	assign leaf[634] = f[407] && !f[359] && f[512] && !f[655];
	assign leaf[635] = f[407] && !f[359] && f[512] && f[655];
	assign leaf[636] = f[407] && f[359] && !f[245] && !f[453];
	assign leaf[637] = f[407] && f[359] && !f[245] && f[453];
	assign leaf[638] = f[407] && f[359] && f[245] && !f[468];
	assign leaf[639] = f[407] && f[359] && f[245] && f[468];
	
	// Tree 41, Classifier 1, Iteration: 4
	assign leaf[640] = !f[437] && !f[346] && !f[578] && !f[300];
	assign leaf[641] = !f[437] && !f[346] && !f[578] && f[300];
	assign leaf[642] = !f[437] && !f[346] && f[578] && !f[293];
	assign leaf[643] = !f[437] && !f[346] && f[578] && f[293];
	assign leaf[644] = !f[437] && f[346] && !f[294] && !f[120];
	assign leaf[645] = !f[437] && f[346] && !f[294] && f[120];
	assign leaf[646] = !f[437] && f[346] && f[294] && !f[435];
	assign leaf[647] = !f[437] && f[346] && f[294] && f[435];
	assign leaf[648] = f[437] && !f[438] && !f[323] && !f[436];
	assign leaf[649] = f[437] && !f[438] && !f[323] && f[436];
	assign leaf[650] = f[437] && !f[438] && f[323] && !f[489];
	assign leaf[651] = f[437] && !f[438] && f[323] && f[489];
	assign leaf[652] = f[437] && f[438] && !f[69];
	assign leaf[653] = f[437] && f[438] && f[69] && !f[383];
	assign leaf[654] = f[437] && f[438] && f[69] && f[383];
	
	// Tree 42, Classifier 2, Iteration: 4
	assign leaf[655] = !f[345] && !f[348] && !f[153] && !f[538];
	assign leaf[656] = !f[345] && !f[348] && !f[153] && f[538];
	assign leaf[657] = !f[345] && !f[348] && f[153] && !f[516];
	assign leaf[658] = !f[345] && !f[348] && f[153] && f[516];
	assign leaf[659] = !f[345] && f[348] && !f[473] && !f[554];
	assign leaf[660] = !f[345] && f[348] && !f[473] && f[554];
	assign leaf[661] = !f[345] && f[348] && f[473] && !f[528];
	assign leaf[662] = !f[345] && f[348] && f[473] && f[528];
	assign leaf[663] = f[345] && !f[583] && !f[501] && !f[568];
	assign leaf[664] = f[345] && !f[583] && !f[501] && f[568];
	assign leaf[665] = f[345] && !f[583] && f[501] && !f[267];
	assign leaf[666] = f[345] && !f[583] && f[501] && f[267];
	assign leaf[667] = f[345] && f[583] && !f[518] && !f[490];
	assign leaf[668] = f[345] && f[583] && !f[518] && f[490];
	assign leaf[669] = f[345] && f[583] && f[518] && !f[430];
	assign leaf[670] = f[345] && f[583] && f[518] && f[430];
	
	// Tree 43, Classifier 3, Iteration: 4
	assign leaf[671] = !f[518] && !f[316] && !f[291] && !f[515];
	assign leaf[672] = !f[518] && !f[316] && !f[291] && f[515];
	assign leaf[673] = !f[518] && !f[316] && f[291] && !f[176];
	assign leaf[674] = !f[518] && !f[316] && f[291] && f[176];
	assign leaf[675] = !f[518] && f[316] && !f[399] && !f[292];
	assign leaf[676] = !f[518] && f[316] && !f[399] && f[292];
	assign leaf[677] = !f[518] && f[316] && f[399] && !f[121];
	assign leaf[678] = !f[518] && f[316] && f[399] && f[121];
	assign leaf[679] = f[518] && !f[624] && !f[463] && !f[352];
	assign leaf[680] = f[518] && !f[624] && !f[463] && f[352];
	assign leaf[681] = f[518] && !f[624] && f[463] && !f[650];
	assign leaf[682] = f[518] && !f[624] && f[463] && f[650];
	assign leaf[683] = f[518] && f[624] && !f[351] && !f[203];
	assign leaf[684] = f[518] && f[624] && !f[351] && f[203];
	assign leaf[685] = f[518] && f[624] && f[351] && !f[485];
	assign leaf[686] = f[518] && f[624] && f[351] && f[485];
	
	// Tree 44, Classifier 4, Iteration: 4
	assign leaf[687] = !f[597] && !f[210] && !f[543] && !f[266];
	assign leaf[688] = !f[597] && !f[210] && !f[543] && f[266];
	assign leaf[689] = !f[597] && !f[210] && f[543] && !f[189];
	assign leaf[690] = !f[597] && !f[210] && f[543] && f[189];
	assign leaf[691] = !f[597] && f[210] && !f[319] && !f[208];
	assign leaf[692] = !f[597] && f[210] && !f[319] && f[208];
	assign leaf[693] = !f[597] && f[210] && f[319] && !f[455];
	assign leaf[694] = !f[597] && f[210] && f[319] && f[455];
	assign leaf[695] = f[597] && !f[163] && !f[220] && !f[156];
	assign leaf[696] = f[597] && !f[163] && !f[220] && f[156];
	assign leaf[697] = f[597] && !f[163] && f[220] && !f[243];
	assign leaf[698] = f[597] && !f[163] && f[220] && f[243];
	assign leaf[699] = f[597] && f[163] && !f[187] && !f[567];
	assign leaf[700] = f[597] && f[163] && !f[187] && f[567];
	assign leaf[701] = f[597] && f[163] && f[187] && !f[213];
	assign leaf[702] = f[597] && f[163] && f[187] && f[213];
	
	// Tree 45, Classifier 5, Iteration: 4
	assign leaf[703] = !f[375] && !f[320] && !f[191] && !f[248];
	assign leaf[704] = !f[375] && !f[320] && !f[191] && f[248];
	assign leaf[705] = !f[375] && !f[320] && f[191] && !f[300];
	assign leaf[706] = !f[375] && !f[320] && f[191] && f[300];
	assign leaf[707] = !f[375] && f[320] && !f[434] && !f[267];
	assign leaf[708] = !f[375] && f[320] && !f[434] && f[267];
	assign leaf[709] = !f[375] && f[320] && f[434] && !f[380];
	assign leaf[710] = !f[375] && f[320] && f[434] && f[380];
	assign leaf[711] = f[375] && !f[486] && !f[297] && !f[299];
	assign leaf[712] = f[375] && !f[486] && !f[297] && f[299];
	assign leaf[713] = f[375] && !f[486] && f[297] && !f[274];
	assign leaf[714] = f[375] && !f[486] && f[297] && f[274];
	assign leaf[715] = f[375] && f[486] && !f[514] && !f[484];
	assign leaf[716] = f[375] && f[486] && !f[514] && f[484];
	assign leaf[717] = f[375] && f[486] && f[514] && !f[458];
	assign leaf[718] = f[375] && f[486] && f[514] && f[458];
	
	// Tree 46, Classifier 6, Iteration: 4
	assign leaf[719] = !f[514] && !f[512] && !f[515] && !f[387];
	assign leaf[720] = !f[514] && !f[512] && !f[515] && f[387];
	assign leaf[721] = !f[514] && !f[512] && f[515] && !f[431];
	assign leaf[722] = !f[514] && !f[512] && f[515] && f[431];
	assign leaf[723] = !f[514] && f[512] && !f[243] && !f[269];
	assign leaf[724] = !f[514] && f[512] && !f[243] && f[269];
	assign leaf[725] = !f[514] && f[512] && f[243] && !f[135];
	assign leaf[726] = !f[514] && f[512] && f[243] && f[135];
	assign leaf[727] = f[514] && !f[270] && !f[272] && !f[296];
	assign leaf[728] = f[514] && !f[270] && !f[272] && f[296];
	assign leaf[729] = f[514] && !f[270] && f[272] && !f[388];
	assign leaf[730] = f[514] && !f[270] && f[272] && f[388];
	assign leaf[731] = f[514] && f[270] && !f[386] && !f[106];
	assign leaf[732] = f[514] && f[270] && !f[386] && f[106];
	assign leaf[733] = f[514] && f[270] && f[386] && !f[241];
	assign leaf[734] = f[514] && f[270] && f[386] && f[241];
	
	// Tree 47, Classifier 7, Iteration: 4
	assign leaf[735] = !f[404] && !f[155] && !f[428] && !f[377];
	assign leaf[736] = !f[404] && !f[155] && !f[428] && f[377];
	assign leaf[737] = !f[404] && !f[155] && f[428] && !f[487];
	assign leaf[738] = !f[404] && !f[155] && f[428] && f[487];
	assign leaf[739] = !f[404] && f[155] && !f[678] && !f[127];
	assign leaf[740] = !f[404] && f[155] && !f[678] && f[127];
	assign leaf[741] = !f[404] && f[155] && f[678] && !f[603];
	assign leaf[742] = !f[404] && f[155] && f[678] && f[603];
	assign leaf[743] = f[404] && !f[412] && !f[441] && !f[345];
	assign leaf[744] = f[404] && !f[412] && !f[441] && f[345];
	assign leaf[745] = f[404] && !f[412] && f[441] && !f[714];
	assign leaf[746] = f[404] && !f[412] && f[441] && f[714];
	assign leaf[747] = f[404] && f[412] && !f[715] && !f[710];
	assign leaf[748] = f[404] && f[412] && !f[715] && f[710];
	assign leaf[749] = f[404] && f[412] && f[715] && !f[322];
	assign leaf[750] = f[404] && f[412] && f[715] && f[322];
	
	// Tree 48, Classifier 8, Iteration: 4
	assign leaf[751] = !f[433] && !f[431] && !f[434] && !f[429];
	assign leaf[752] = !f[433] && !f[431] && !f[434] && f[429];
	assign leaf[753] = !f[433] && !f[431] && f[434] && !f[377];
	assign leaf[754] = !f[433] && !f[431] && f[434] && f[377];
	assign leaf[755] = !f[433] && f[431] && !f[658] && !f[655];
	assign leaf[756] = !f[433] && f[431] && !f[658] && f[655];
	assign leaf[757] = !f[433] && f[431] && f[658] && !f[374];
	assign leaf[758] = !f[433] && f[431] && f[658] && f[374];
	assign leaf[759] = f[433] && !f[657] && !f[303] && !f[629];
	assign leaf[760] = f[433] && !f[657] && !f[303] && f[629];
	assign leaf[761] = f[433] && !f[657] && f[303] && !f[408];
	assign leaf[762] = f[433] && !f[657] && f[303] && f[408];
	assign leaf[763] = f[433] && f[657] && !f[515] && !f[512];
	assign leaf[764] = f[433] && f[657] && !f[515] && f[512];
	assign leaf[765] = f[433] && f[657] && f[515] && !f[290];
	assign leaf[766] = f[433] && f[657] && f[515] && f[290];
	
	// Tree 49, Classifier 9, Iteration: 4
	assign leaf[767] = !f[598] && !f[372] && !f[398] && !f[346];
	assign leaf[768] = !f[598] && !f[372] && !f[398] && f[346];
	assign leaf[769] = !f[598] && !f[372] && f[398] && !f[209];
	assign leaf[770] = !f[598] && !f[372] && f[398] && f[209];
	assign leaf[771] = !f[598] && f[372] && !f[210] && !f[238];
	assign leaf[772] = !f[598] && f[372] && !f[210] && f[238];
	assign leaf[773] = !f[598] && f[372] && f[210] && !f[347];
	assign leaf[774] = !f[598] && f[372] && f[210] && f[347];
	assign leaf[775] = f[598] && !f[708] && !f[706] && !f[709];
	assign leaf[776] = f[598] && !f[708] && !f[706] && f[709];
	assign leaf[777] = f[598] && !f[708] && f[706] && !f[406];
	assign leaf[778] = f[598] && !f[708] && f[706] && f[406];
	assign leaf[779] = f[598] && f[708] && !f[405] && !f[350];
	assign leaf[780] = f[598] && f[708] && !f[405] && f[350];
	assign leaf[781] = f[598] && f[708] && f[405] && !f[233];
	assign leaf[782] = f[598] && f[708] && f[405] && f[233];
	
	// Tree 50, Classifier 0, Iteration: 5
	assign leaf[783] = !f[435] && !f[379] && !f[598] && !f[539];
	assign leaf[784] = !f[435] && !f[379] && !f[598] && f[539];
	assign leaf[785] = !f[435] && !f[379] && f[598] && !f[489];
	assign leaf[786] = !f[435] && !f[379] && f[598] && f[489];
	assign leaf[787] = !f[435] && f[379] && !f[331] && !f[329];
	assign leaf[788] = !f[435] && f[379] && !f[331] && f[329];
	assign leaf[789] = !f[435] && f[379] && f[331] && !f[265];
	assign leaf[790] = !f[435] && f[379] && f[331] && f[265];
	assign leaf[791] = f[435] && !f[386] && !f[540] && !f[539];
	assign leaf[792] = f[435] && !f[386] && !f[540] && f[539];
	assign leaf[793] = f[435] && !f[386] && f[540] && !f[434];
	assign leaf[794] = f[435] && !f[386] && f[540] && f[434];
	assign leaf[795] = f[435] && f[386] && !f[322] && !f[625];
	assign leaf[796] = f[435] && f[386] && !f[322] && f[625];
	assign leaf[797] = f[435] && f[386] && f[322] && !f[433];
	assign leaf[798] = f[435] && f[386] && f[322] && f[433];
	
	// Tree 51, Classifier 1, Iteration: 5
	assign leaf[799] = !f[382] && !f[465] && !f[378] && !f[379];
	assign leaf[800] = !f[382] && !f[465] && !f[378] && f[379];
	assign leaf[801] = !f[382] && !f[465] && f[378] && !f[206];
	assign leaf[802] = !f[382] && !f[465] && f[378] && f[206];
	assign leaf[803] = !f[382] && f[465] && !f[466] && !f[518];
	assign leaf[804] = !f[382] && f[465] && !f[466] && f[518];
	assign leaf[805] = !f[382] && f[465] && f[466] && !f[98];
	assign leaf[806] = !f[382] && f[465] && f[466] && f[98];
	assign leaf[807] = f[382] && !f[162] && !f[355] && !f[488];
	assign leaf[808] = f[382] && !f[162] && !f[355] && f[488];
	assign leaf[809] = f[382] && !f[162] && f[355];
	assign leaf[810] = f[382] && f[162] && !f[269] && !f[296];
	assign leaf[811] = f[382] && f[162] && !f[269] && f[296];
	assign leaf[812] = f[382] && f[162] && f[269] && !f[320];
	assign leaf[813] = f[382] && f[162] && f[269] && f[320];
	
	// Tree 52, Classifier 2, Iteration: 5
	assign leaf[814] = !f[543] && !f[512] && !f[99] && !f[514];
	assign leaf[815] = !f[543] && !f[512] && !f[99] && f[514];
	assign leaf[816] = !f[543] && !f[512] && f[99] && !f[351];
	assign leaf[817] = !f[543] && !f[512] && f[99] && f[351];
	assign leaf[818] = !f[543] && f[512] && !f[319] && !f[316];
	assign leaf[819] = !f[543] && f[512] && !f[319] && f[316];
	assign leaf[820] = !f[543] && f[512] && f[319] && !f[630];
	assign leaf[821] = !f[543] && f[512] && f[319] && f[630];
	assign leaf[822] = f[543] && !f[346] && !f[181] && !f[126];
	assign leaf[823] = f[543] && !f[346] && !f[181] && f[126];
	assign leaf[824] = f[543] && !f[346] && f[181] && !f[371];
	assign leaf[825] = f[543] && !f[346] && f[181] && f[371];
	assign leaf[826] = f[543] && f[346] && !f[318] && !f[426];
	assign leaf[827] = f[543] && f[346] && !f[318] && f[426];
	assign leaf[828] = f[543] && f[346] && f[318] && !f[374];
	assign leaf[829] = f[543] && f[346] && f[318] && f[374];
	
	// Tree 53, Classifier 3, Iteration: 5
	assign leaf[830] = !f[152] && !f[180] && !f[563] && !f[507];
	assign leaf[831] = !f[152] && !f[180] && !f[563] && f[507];
	assign leaf[832] = !f[152] && !f[180] && f[563] && !f[482];
	assign leaf[833] = !f[152] && !f[180] && f[563] && f[482];
	assign leaf[834] = !f[152] && f[180] && !f[317] && !f[515];
	assign leaf[835] = !f[152] && f[180] && !f[317] && f[515];
	assign leaf[836] = !f[152] && f[180] && f[317] && !f[228];
	assign leaf[837] = !f[152] && f[180] && f[317] && f[228];
	assign leaf[838] = f[152] && !f[485] && !f[296] && !f[239];
	assign leaf[839] = f[152] && !f[485] && !f[296] && f[239];
	assign leaf[840] = f[152] && !f[485] && f[296] && !f[516];
	assign leaf[841] = f[152] && !f[485] && f[296] && f[516];
	assign leaf[842] = f[152] && f[485] && !f[295] && !f[678];
	assign leaf[843] = f[152] && f[485] && !f[295] && f[678];
	assign leaf[844] = f[152] && f[485] && f[295] && !f[431];
	assign leaf[845] = f[152] && f[485] && f[295] && f[431];
	
	// Tree 54, Classifier 4, Iteration: 5
	assign leaf[846] = !f[464] && !f[183] && !f[436] && !f[295];
	assign leaf[847] = !f[464] && !f[183] && !f[436] && f[295];
	assign leaf[848] = !f[464] && !f[183] && f[436] && !f[575];
	assign leaf[849] = !f[464] && !f[183] && f[436] && f[575];
	assign leaf[850] = !f[464] && f[183] && !f[185] && !f[246];
	assign leaf[851] = !f[464] && f[183] && !f[185] && f[246];
	assign leaf[852] = !f[464] && f[183] && f[185] && !f[368];
	assign leaf[853] = !f[464] && f[183] && f[185] && f[368];
	assign leaf[854] = f[464] && !f[210] && !f[154] && !f[266];
	assign leaf[855] = f[464] && !f[210] && !f[154] && f[266];
	assign leaf[856] = f[464] && !f[210] && f[154] && !f[155];
	assign leaf[857] = f[464] && !f[210] && f[154] && f[155];
	assign leaf[858] = f[464] && f[210] && !f[213] && !f[292];
	assign leaf[859] = f[464] && f[210] && !f[213] && f[292];
	assign leaf[860] = f[464] && f[210] && f[213] && !f[442];
	assign leaf[861] = f[464] && f[210] && f[213] && f[442];
	
	// Tree 55, Classifier 5, Iteration: 5
	assign leaf[862] = !f[327] && !f[296] && !f[517] && !f[330];
	assign leaf[863] = !f[327] && !f[296] && !f[517] && f[330];
	assign leaf[864] = !f[327] && !f[296] && f[517] && !f[217];
	assign leaf[865] = !f[327] && !f[296] && f[517] && f[217];
	assign leaf[866] = !f[327] && f[296] && !f[273] && !f[218];
	assign leaf[867] = !f[327] && f[296] && !f[273] && f[218];
	assign leaf[868] = !f[327] && f[296] && f[273] && !f[358];
	assign leaf[869] = !f[327] && f[296] && f[273] && f[358];
	assign leaf[870] = f[327] && !f[323] && !f[305] && !f[382];
	assign leaf[871] = f[327] && !f[323] && !f[305] && f[382];
	assign leaf[872] = f[327] && !f[323] && f[305] && !f[381];
	assign leaf[873] = f[327] && !f[323] && f[305] && f[381];
	assign leaf[874] = f[327] && f[323] && !f[409] && !f[522];
	assign leaf[875] = f[327] && f[323] && !f[409] && f[522];
	assign leaf[876] = f[327] && f[323] && f[409] && !f[248];
	assign leaf[877] = f[327] && f[323] && f[409] && f[248];
	
	// Tree 56, Classifier 6, Iteration: 5
	assign leaf[878] = !f[270] && !f[543] && !f[541] && !f[516];
	assign leaf[879] = !f[270] && !f[543] && !f[541] && f[516];
	assign leaf[880] = !f[270] && !f[543] && f[541] && !f[244];
	assign leaf[881] = !f[270] && !f[543] && f[541] && f[244];
	assign leaf[882] = !f[270] && f[543] && !f[574] && !f[601];
	assign leaf[883] = !f[270] && f[543] && !f[574] && f[601];
	assign leaf[884] = !f[270] && f[543] && f[574] && !f[245];
	assign leaf[885] = !f[270] && f[543] && f[574] && f[245];
	assign leaf[886] = f[270] && !f[92] && !f[136] && !f[94];
	assign leaf[887] = f[270] && !f[92] && !f[136] && f[94];
	assign leaf[888] = f[270] && !f[92] && f[136] && !f[429];
	assign leaf[889] = f[270] && !f[92] && f[136] && f[429];
	assign leaf[890] = f[270] && f[92] && !f[123] && !f[150];
	assign leaf[891] = f[270] && f[92] && !f[123] && f[150];
	assign leaf[892] = f[270] && f[92] && f[123];
	
	// Tree 57, Classifier 7, Iteration: 5
	assign leaf[893] = !f[404] && !f[157] && !f[269] && !f[461];
	assign leaf[894] = !f[404] && !f[157] && !f[269] && f[461];
	assign leaf[895] = !f[404] && !f[157] && f[269] && !f[541];
	assign leaf[896] = !f[404] && !f[157] && f[269] && f[541];
	assign leaf[897] = !f[404] && f[157] && !f[203] && !f[679];
	assign leaf[898] = !f[404] && f[157] && !f[203] && f[679];
	assign leaf[899] = !f[404] && f[157] && f[203] && !f[606];
	assign leaf[900] = !f[404] && f[157] && f[203] && f[606];
	assign leaf[901] = f[404] && !f[155] && !f[412] && !f[296];
	assign leaf[902] = f[404] && !f[155] && !f[412] && f[296];
	assign leaf[903] = f[404] && !f[155] && f[412] && !f[323];
	assign leaf[904] = f[404] && !f[155] && f[412] && f[323];
	assign leaf[905] = f[404] && f[155];
	
	// Tree 58, Classifier 8, Iteration: 5
	assign leaf[906] = !f[433] && !f[431] && !f[378] && !f[405];
	assign leaf[907] = !f[433] && !f[431] && !f[378] && f[405];
	assign leaf[908] = !f[433] && !f[431] && f[378] && !f[489];
	assign leaf[909] = !f[433] && !f[431] && f[378] && f[489];
	assign leaf[910] = !f[433] && f[431] && !f[548] && !f[400];
	assign leaf[911] = !f[433] && f[431] && !f[548] && f[400];
	assign leaf[912] = !f[433] && f[431] && f[548] && !f[434];
	assign leaf[913] = !f[433] && f[431] && f[548] && f[434];
	assign leaf[914] = f[433] && !f[348] && !f[375] && !f[321];
	assign leaf[915] = f[433] && !f[348] && !f[375] && f[321];
	assign leaf[916] = f[433] && !f[348] && f[375] && !f[429];
	assign leaf[917] = f[433] && !f[348] && f[375] && f[429];
	assign leaf[918] = f[433] && f[348] && !f[402] && !f[294];
	assign leaf[919] = f[433] && f[348] && !f[402] && f[294];
	assign leaf[920] = f[433] && f[348] && f[402] && !f[289];
	assign leaf[921] = f[433] && f[348] && f[402] && f[289];
	
	// Tree 59, Classifier 9, Iteration: 5
	assign leaf[922] = !f[570] && !f[624] && !f[212] && !f[692];
	assign leaf[923] = !f[570] && !f[624] && !f[212] && f[692];
	assign leaf[924] = !f[570] && !f[624] && f[212] && !f[205];
	assign leaf[925] = !f[570] && !f[624] && f[212] && f[205];
	assign leaf[926] = !f[570] && f[624] && !f[706] && !f[238];
	assign leaf[927] = !f[570] && f[624] && !f[706] && f[238];
	assign leaf[928] = !f[570] && f[624] && f[706];
	assign leaf[929] = f[570] && !f[680] && !f[719] && !f[340];
	assign leaf[930] = f[570] && !f[680] && !f[719] && f[340];
	assign leaf[931] = f[570] && !f[680] && f[719] && !f[573];
	assign leaf[932] = f[570] && !f[680] && f[719] && f[573];
	assign leaf[933] = f[570] && f[680] && !f[374] && !f[348];
	assign leaf[934] = f[570] && f[680] && !f[374] && f[348];
	assign leaf[935] = f[570] && f[680] && f[374] && !f[214];
	assign leaf[936] = f[570] && f[680] && f[374] && f[214];
	
	// Tree 60, Classifier 0, Iteration: 6
	assign leaf[937] = !f[434] && !f[455] && !f[457] && !f[425];
	assign leaf[938] = !f[434] && !f[455] && !f[457] && f[425];
	assign leaf[939] = !f[434] && !f[455] && f[457] && !f[628];
	assign leaf[940] = !f[434] && !f[455] && f[457] && f[628];
	assign leaf[941] = !f[434] && f[455] && !f[626] && !f[410];
	assign leaf[942] = !f[434] && f[455] && !f[626] && f[410];
	assign leaf[943] = !f[434] && f[455] && f[626] && !f[378];
	assign leaf[944] = !f[434] && f[455] && f[626] && f[378];
	assign leaf[945] = f[434] && !f[385] && !f[359];
	assign leaf[946] = f[434] && !f[385] && f[359] && !f[185];
	assign leaf[947] = f[434] && !f[385] && f[359] && f[185];
	assign leaf[948] = f[434] && f[385] && !f[409] && !f[655];
	assign leaf[949] = f[434] && f[385] && !f[409] && f[655];
	assign leaf[950] = f[434] && f[385] && f[409] && !f[274];
	assign leaf[951] = f[434] && f[385] && f[409] && f[274];
	
	// Tree 61, Classifier 1, Iteration: 6
	assign leaf[952] = !f[323] && !f[322] && !f[211] && !f[650];
	assign leaf[953] = !f[323] && !f[322] && !f[211] && f[650];
	assign leaf[954] = !f[323] && !f[322] && f[211] && !f[378];
	assign leaf[955] = !f[323] && !f[322] && f[211] && f[378];
	assign leaf[956] = !f[323] && f[322] && !f[627] && !f[380];
	assign leaf[957] = !f[323] && f[322] && !f[627] && f[380];
	assign leaf[958] = !f[323] && f[322] && f[627] && !f[126];
	assign leaf[959] = !f[323] && f[322] && f[627] && f[126];
	assign leaf[960] = f[323] && !f[494] && !f[234] && !f[402];
	assign leaf[961] = f[323] && !f[494] && !f[234] && f[402];
	assign leaf[962] = f[323] && !f[494] && f[234] && !f[324];
	assign leaf[963] = f[323] && !f[494] && f[234] && f[324];
	assign leaf[964] = f[323] && f[494] && !f[71] && !f[98];
	assign leaf[965] = f[323] && f[494] && !f[71] && f[98];
	assign leaf[966] = f[323] && f[494] && f[71];
	
	// Tree 62, Classifier 2, Iteration: 6
	assign leaf[967] = !f[346] && !f[543] && !f[485] && !f[514];
	assign leaf[968] = !f[346] && !f[543] && !f[485] && f[514];
	assign leaf[969] = !f[346] && !f[543] && f[485] && !f[343];
	assign leaf[970] = !f[346] && !f[543] && f[485] && f[343];
	assign leaf[971] = !f[346] && f[543] && !f[154] && !f[653];
	assign leaf[972] = !f[346] && f[543] && !f[154] && f[653];
	assign leaf[973] = !f[346] && f[543] && f[154] && !f[320];
	assign leaf[974] = !f[346] && f[543] && f[154] && f[320];
	assign leaf[975] = f[346] && !f[582] && !f[527] && !f[637];
	assign leaf[976] = f[346] && !f[582] && !f[527] && f[637];
	assign leaf[977] = f[346] && !f[582] && f[527] && !f[604];
	assign leaf[978] = f[346] && !f[582] && f[527] && f[604];
	assign leaf[979] = f[346] && f[582] && !f[633] && !f[522];
	assign leaf[980] = f[346] && f[582] && !f[633] && f[522];
	assign leaf[981] = f[346] && f[582] && f[633] && !f[547];
	assign leaf[982] = f[346] && f[582] && f[633] && f[547];
	
	// Tree 63, Classifier 3, Iteration: 6
	assign leaf[983] = !f[490] && !f[343] && !f[485] && !f[263];
	assign leaf[984] = !f[490] && !f[343] && !f[485] && f[263];
	assign leaf[985] = !f[490] && !f[343] && f[485] && !f[203];
	assign leaf[986] = !f[490] && !f[343] && f[485] && f[203];
	assign leaf[987] = !f[490] && f[343] && !f[287] && !f[149];
	assign leaf[988] = !f[490] && f[343] && !f[287] && f[149];
	assign leaf[989] = !f[490] && f[343] && f[287] && !f[289];
	assign leaf[990] = !f[490] && f[343] && f[287] && f[289];
	assign leaf[991] = f[490] && !f[324] && !f[682] && !f[203];
	assign leaf[992] = f[490] && !f[324] && !f[682] && f[203];
	assign leaf[993] = f[490] && !f[324] && f[682] && !f[545];
	assign leaf[994] = f[490] && !f[324] && f[682] && f[545];
	assign leaf[995] = f[490] && f[324] && !f[181] && !f[101];
	assign leaf[996] = f[490] && f[324] && !f[181] && f[101];
	assign leaf[997] = f[490] && f[324] && f[181] && !f[654];
	assign leaf[998] = f[490] && f[324] && f[181] && f[654];
	
	// Tree 64, Classifier 4, Iteration: 6
	assign leaf[999] = !f[569] && !f[427] && !f[374] && !f[373];
	assign leaf[1000] = !f[569] && !f[427] && !f[374] && f[373];
	assign leaf[1001] = !f[569] && !f[427] && f[374] && !f[551];
	assign leaf[1002] = !f[569] && !f[427] && f[374] && f[551];
	assign leaf[1003] = !f[569] && f[427] && !f[374] && !f[238];
	assign leaf[1004] = !f[569] && f[427] && !f[374] && f[238];
	assign leaf[1005] = !f[569] && f[427] && f[374] && !f[623];
	assign leaf[1006] = !f[569] && f[427] && f[374] && f[623];
	assign leaf[1007] = f[569] && !f[163] && !f[600] && !f[400];
	assign leaf[1008] = f[569] && !f[163] && !f[600] && f[400];
	assign leaf[1009] = f[569] && !f[163] && f[600] && !f[710];
	assign leaf[1010] = f[569] && !f[163] && f[600] && f[710];
	assign leaf[1011] = f[569] && f[163] && !f[595] && !f[213];
	assign leaf[1012] = f[569] && f[163] && !f[595] && f[213];
	assign leaf[1013] = f[569] && f[163] && f[595] && !f[567];
	assign leaf[1014] = f[569] && f[163] && f[595] && f[567];
	
	// Tree 65, Classifier 5, Iteration: 6
	assign leaf[1015] = !f[489] && !f[298] && !f[267] && !f[301];
	assign leaf[1016] = !f[489] && !f[298] && !f[267] && f[301];
	assign leaf[1017] = !f[489] && !f[298] && f[267] && !f[243];
	assign leaf[1018] = !f[489] && !f[298] && f[267] && f[243];
	assign leaf[1019] = !f[489] && f[298] && !f[275] && !f[304];
	assign leaf[1020] = !f[489] && f[298] && !f[275] && f[304];
	assign leaf[1021] = !f[489] && f[298] && f[275] && !f[186];
	assign leaf[1022] = !f[489] && f[298] && f[275] && f[186];
	assign leaf[1023] = f[489] && !f[380] && !f[410] && !f[378];
	assign leaf[1024] = f[489] && !f[380] && !f[410] && f[378];
	assign leaf[1025] = f[489] && !f[380] && f[410] && !f[352];
	assign leaf[1026] = f[489] && !f[380] && f[410] && f[352];
	assign leaf[1027] = f[489] && f[380] && !f[510] && !f[537];
	assign leaf[1028] = f[489] && f[380] && !f[510] && f[537];
	assign leaf[1029] = f[489] && f[380] && f[510] && !f[461];
	assign leaf[1030] = f[489] && f[380] && f[510] && f[461];
	
	// Tree 66, Classifier 6, Iteration: 6
	assign leaf[1031] = !f[270] && !f[486] && !f[484] && !f[487];
	assign leaf[1032] = !f[270] && !f[486] && !f[484] && f[487];
	assign leaf[1033] = !f[270] && !f[486] && f[484] && !f[244];
	assign leaf[1034] = !f[270] && !f[486] && f[484] && f[244];
	assign leaf[1035] = !f[270] && f[486] && !f[272] && !f[296];
	assign leaf[1036] = !f[270] && f[486] && !f[272] && f[296];
	assign leaf[1037] = !f[270] && f[486] && f[272] && !f[359];
	assign leaf[1038] = !f[270] && f[486] && f[272] && f[359];
	assign leaf[1039] = f[270] && !f[386] && !f[107] && !f[359];
	assign leaf[1040] = f[270] && !f[386] && !f[107] && f[359];
	assign leaf[1041] = f[270] && !f[386] && f[107];
	assign leaf[1042] = f[270] && f[386] && !f[122] && !f[119];
	assign leaf[1043] = f[270] && f[386] && !f[122] && f[119];
	assign leaf[1044] = f[270] && f[386] && f[122] && !f[212];
	assign leaf[1045] = f[270] && f[386] && f[122] && f[212];
	
	// Tree 67, Classifier 7, Iteration: 6
	assign leaf[1046] = !f[377] && !f[459] && !f[512] && !f[158];
	assign leaf[1047] = !f[377] && !f[459] && !f[512] && f[158];
	assign leaf[1048] = !f[377] && !f[459] && f[512] && !f[715];
	assign leaf[1049] = !f[377] && !f[459] && f[512] && f[715];
	assign leaf[1050] = !f[377] && f[459] && !f[373] && !f[324];
	assign leaf[1051] = !f[377] && f[459] && !f[373] && f[324];
	assign leaf[1052] = !f[377] && f[459] && f[373] && !f[285];
	assign leaf[1053] = !f[377] && f[459] && f[373] && f[285];
	assign leaf[1054] = f[377] && !f[339] && !f[385] && !f[517];
	assign leaf[1055] = f[377] && !f[339] && !f[385] && f[517];
	assign leaf[1056] = f[377] && !f[339] && f[385] && !f[186];
	assign leaf[1057] = f[377] && !f[339] && f[385] && f[186];
	assign leaf[1058] = f[377] && f[339] && !f[257] && !f[269];
	assign leaf[1059] = f[377] && f[339] && !f[257] && f[269];
	assign leaf[1060] = f[377] && f[339] && f[257];
	
	// Tree 68, Classifier 8, Iteration: 6
	assign leaf[1061] = !f[406] && !f[404] && !f[430] && !f[350];
	assign leaf[1062] = !f[406] && !f[404] && !f[430] && f[350];
	assign leaf[1063] = !f[406] && !f[404] && f[430] && !f[493];
	assign leaf[1064] = !f[406] && !f[404] && f[430] && f[493];
	assign leaf[1065] = !f[406] && f[404] && !f[408] && !f[522];
	assign leaf[1066] = !f[406] && f[404] && !f[408] && f[522];
	assign leaf[1067] = !f[406] && f[404] && f[408] && !f[656];
	assign leaf[1068] = !f[406] && f[404] && f[408] && f[656];
	assign leaf[1069] = f[406] && !f[487] && !f[485] && !f[516];
	assign leaf[1070] = f[406] && !f[487] && !f[485] && f[516];
	assign leaf[1071] = f[406] && !f[487] && f[485] && !f[437];
	assign leaf[1072] = f[406] && !f[487] && f[485] && f[437];
	assign leaf[1073] = f[406] && f[487] && !f[428] && !f[348];
	assign leaf[1074] = f[406] && f[487] && !f[428] && f[348];
	assign leaf[1075] = f[406] && f[487] && f[428] && !f[625];
	assign leaf[1076] = f[406] && f[487] && f[428] && f[625];
	
	// Tree 69, Classifier 9, Iteration: 6
	assign leaf[1077] = !f[569] && !f[354] && !f[157] && !f[290];
	assign leaf[1078] = !f[569] && !f[354] && !f[157] && f[290];
	assign leaf[1079] = !f[569] && !f[354] && f[157] && !f[384];
	assign leaf[1080] = !f[569] && !f[354] && f[157] && f[384];
	assign leaf[1081] = !f[569] && f[354] && !f[406] && !f[487];
	assign leaf[1082] = !f[569] && f[354] && !f[406] && f[487];
	assign leaf[1083] = !f[569] && f[354] && f[406] && !f[623];
	assign leaf[1084] = !f[569] && f[354] && f[406] && f[623];
	assign leaf[1085] = f[569] && !f[368] && !f[706] && !f[689];
	assign leaf[1086] = f[569] && !f[368] && !f[706] && f[689];
	assign leaf[1087] = f[569] && !f[368] && f[706] && !f[376];
	assign leaf[1088] = f[569] && !f[368] && f[706] && f[376];
	assign leaf[1089] = f[569] && f[368] && !f[355];
	assign leaf[1090] = f[569] && f[368] && f[355] && !f[340];
	assign leaf[1091] = f[569] && f[368] && f[355] && f[340];
	
	// Tree 70, Classifier 0, Iteration: 7
	assign leaf[1092] = !f[408] && !f[461] && !f[352] && !f[214];
	assign leaf[1093] = !f[408] && !f[461] && !f[352] && f[214];
	assign leaf[1094] = !f[408] && !f[461] && f[352] && !f[265];
	assign leaf[1095] = !f[408] && !f[461] && f[352] && f[265];
	assign leaf[1096] = !f[408] && f[461] && !f[386] && !f[657];
	assign leaf[1097] = !f[408] && f[461] && !f[386] && f[657];
	assign leaf[1098] = !f[408] && f[461] && f[386] && !f[293];
	assign leaf[1099] = !f[408] && f[461] && f[386] && f[293];
	assign leaf[1100] = f[408] && !f[484] && !f[514] && !f[481];
	assign leaf[1101] = f[408] && !f[484] && !f[514] && f[481];
	assign leaf[1102] = f[408] && !f[484] && f[514] && !f[434];
	assign leaf[1103] = f[408] && !f[484] && f[514] && f[434];
	assign leaf[1104] = f[408] && f[484] && !f[626] && !f[331];
	assign leaf[1105] = f[408] && f[484] && !f[626] && f[331];
	assign leaf[1106] = f[408] && f[484] && f[626] && !f[433];
	assign leaf[1107] = f[408] && f[484] && f[626] && f[433];
	
	// Tree 71, Classifier 1, Iteration: 7
	assign leaf[1108] = !f[323] && !f[212] && !f[322] && !f[650];
	assign leaf[1109] = !f[323] && !f[212] && !f[322] && f[650];
	assign leaf[1110] = !f[323] && !f[212] && f[322] && !f[380];
	assign leaf[1111] = !f[323] && !f[212] && f[322] && f[380];
	assign leaf[1112] = !f[323] && f[212] && !f[406] && !f[620];
	assign leaf[1113] = !f[323] && f[212] && !f[406] && f[620];
	assign leaf[1114] = !f[323] && f[212] && f[406] && !f[437];
	assign leaf[1115] = !f[323] && f[212] && f[406] && f[437];
	assign leaf[1116] = f[323] && !f[430] && !f[434] && !f[349];
	assign leaf[1117] = f[323] && !f[430] && !f[434] && f[349];
	assign leaf[1118] = f[323] && !f[430] && f[434] && !f[205];
	assign leaf[1119] = f[323] && !f[430] && f[434] && f[205];
	assign leaf[1120] = f[323] && f[430] && !f[236] && !f[189];
	assign leaf[1121] = f[323] && f[430] && !f[236] && f[189];
	assign leaf[1122] = f[323] && f[430] && f[236] && !f[347];
	assign leaf[1123] = f[323] && f[430] && f[236] && f[347];
	
	// Tree 72, Classifier 2, Iteration: 7
	assign leaf[1124] = !f[319] && !f[344] && !f[321] && !f[127];
	assign leaf[1125] = !f[319] && !f[344] && !f[321] && f[127];
	assign leaf[1126] = !f[319] && !f[344] && f[321] && !f[499];
	assign leaf[1127] = !f[319] && !f[344] && f[321] && f[499];
	assign leaf[1128] = !f[319] && f[344] && !f[316] && !f[425];
	assign leaf[1129] = !f[319] && f[344] && !f[316] && f[425];
	assign leaf[1130] = !f[319] && f[344] && f[316] && !f[372];
	assign leaf[1131] = !f[319] && f[344] && f[316] && f[372];
	assign leaf[1132] = f[319] && !f[473] && !f[581] && !f[527];
	assign leaf[1133] = f[319] && !f[473] && !f[581] && f[527];
	assign leaf[1134] = f[319] && !f[473] && f[581] && !f[490];
	assign leaf[1135] = f[319] && !f[473] && f[581] && f[490];
	assign leaf[1136] = f[319] && f[473] && !f[454] && !f[539];
	assign leaf[1137] = f[319] && f[473] && !f[454] && f[539];
	assign leaf[1138] = f[319] && f[473] && f[454];
	
	// Tree 73, Classifier 3, Iteration: 7
	assign leaf[1139] = !f[177] && !f[623] && !f[122] && !f[678];
	assign leaf[1140] = !f[177] && !f[623] && !f[122] && f[678];
	assign leaf[1141] = !f[177] && !f[623] && f[122] && !f[629];
	assign leaf[1142] = !f[177] && !f[623] && f[122] && f[629];
	assign leaf[1143] = !f[177] && f[623] && !f[324] && !f[511];
	assign leaf[1144] = !f[177] && f[623] && !f[324] && f[511];
	assign leaf[1145] = !f[177] && f[623] && f[324] && !f[486];
	assign leaf[1146] = !f[177] && f[623] && f[324] && f[486];
	assign leaf[1147] = f[177] && !f[288] && !f[657] && !f[320];
	assign leaf[1148] = f[177] && !f[288] && !f[657] && f[320];
	assign leaf[1149] = f[177] && !f[288] && f[657] && !f[314];
	assign leaf[1150] = f[177] && !f[288] && f[657] && f[314];
	assign leaf[1151] = f[177] && f[288] && !f[264] && !f[344];
	assign leaf[1152] = f[177] && f[288] && !f[264] && f[344];
	assign leaf[1153] = f[177] && f[288] && f[264] && !f[371];
	assign leaf[1154] = f[177] && f[288] && f[264] && f[371];
	
	// Tree 74, Classifier 4, Iteration: 7
	assign leaf[1155] = !f[401] && !f[598] && !f[238] && !f[182];
	assign leaf[1156] = !f[401] && !f[598] && !f[238] && f[182];
	assign leaf[1157] = !f[401] && !f[598] && f[238] && !f[430];
	assign leaf[1158] = !f[401] && !f[598] && f[238] && f[430];
	assign leaf[1159] = !f[401] && f[598] && !f[163] && !f[681];
	assign leaf[1160] = !f[401] && f[598] && !f[163] && f[681];
	assign leaf[1161] = !f[401] && f[598] && f[163] && !f[595];
	assign leaf[1162] = !f[401] && f[598] && f[163] && f[595];
	assign leaf[1163] = f[401] && !f[552] && !f[462] && !f[626];
	assign leaf[1164] = f[401] && !f[552] && !f[462] && f[626];
	assign leaf[1165] = f[401] && !f[552] && f[462] && !f[567];
	assign leaf[1166] = f[401] && !f[552] && f[462] && f[567];
	assign leaf[1167] = f[401] && f[552] && !f[664] && !f[454];
	assign leaf[1168] = f[401] && f[552] && !f[664] && f[454];
	assign leaf[1169] = f[401] && f[552] && f[664] && !f[209];
	assign leaf[1170] = f[401] && f[552] && f[664] && f[209];
	
	// Tree 75, Classifier 5, Iteration: 7
	assign leaf[1171] = !f[490] && !f[297] && !f[300] && !f[186];
	assign leaf[1172] = !f[490] && !f[297] && !f[300] && f[186];
	assign leaf[1173] = !f[490] && !f[297] && f[300] && !f[328];
	assign leaf[1174] = !f[490] && !f[297] && f[300] && f[328];
	assign leaf[1175] = !f[490] && f[297] && !f[294] && !f[277];
	assign leaf[1176] = !f[490] && f[297] && !f[294] && f[277];
	assign leaf[1177] = !f[490] && f[297] && f[294] && !f[241];
	assign leaf[1178] = !f[490] && f[297] && f[294] && f[241];
	assign leaf[1179] = f[490] && !f[381] && !f[245] && !f[379];
	assign leaf[1180] = f[490] && !f[381] && !f[245] && f[379];
	assign leaf[1181] = f[490] && !f[381] && f[245] && !f[384];
	assign leaf[1182] = f[490] && !f[381] && f[245] && f[384];
	assign leaf[1183] = f[490] && f[381] && !f[435] && !f[510];
	assign leaf[1184] = f[490] && f[381] && !f[435] && f[510];
	assign leaf[1185] = f[490] && f[381] && f[435] && !f[221];
	assign leaf[1186] = f[490] && f[381] && f[435] && f[221];
	
	// Tree 76, Classifier 6, Iteration: 7
	assign leaf[1187] = !f[242] && !f[572] && !f[388] && !f[131];
	assign leaf[1188] = !f[242] && !f[572] && !f[388] && f[131];
	assign leaf[1189] = !f[242] && !f[572] && f[388] && !f[329];
	assign leaf[1190] = !f[242] && !f[572] && f[388] && f[329];
	assign leaf[1191] = !f[242] && f[572] && !f[655] && !f[295];
	assign leaf[1192] = !f[242] && f[572] && !f[655] && f[295];
	assign leaf[1193] = !f[242] && f[572] && f[655] && !f[131];
	assign leaf[1194] = !f[242] && f[572] && f[655] && f[131];
	assign leaf[1195] = f[242] && !f[133] && !f[93] && !f[103];
	assign leaf[1196] = f[242] && !f[133] && !f[93] && f[103];
	assign leaf[1197] = f[242] && !f[133] && f[93] && !f[125];
	assign leaf[1198] = f[242] && !f[133] && f[93] && f[125];
	assign leaf[1199] = f[242] && f[133] && !f[298] && !f[513];
	assign leaf[1200] = f[242] && f[133] && !f[298] && f[513];
	assign leaf[1201] = f[242] && f[133] && f[298] && !f[326];
	assign leaf[1202] = f[242] && f[133] && f[298] && f[326];
	
	// Tree 77, Classifier 7, Iteration: 7
	assign leaf[1203] = !f[154] && !f[432] && !f[513] && !f[378];
	assign leaf[1204] = !f[154] && !f[432] && !f[513] && f[378];
	assign leaf[1205] = !f[154] && !f[432] && f[513] && !f[399];
	assign leaf[1206] = !f[154] && !f[432] && f[513] && f[399];
	assign leaf[1207] = !f[154] && f[432] && !f[232] && !f[205];
	assign leaf[1208] = !f[154] && f[432] && !f[232] && f[205];
	assign leaf[1209] = !f[154] && f[432] && f[232] && !f[578];
	assign leaf[1210] = !f[154] && f[432] && f[232] && f[578];
	assign leaf[1211] = f[154] && !f[577] && !f[679] && !f[296];
	assign leaf[1212] = f[154] && !f[577] && !f[679] && f[296];
	assign leaf[1213] = f[154] && !f[577] && f[679] && !f[571];
	assign leaf[1214] = f[154] && !f[577] && f[679] && f[571];
	assign leaf[1215] = f[154] && f[577] && !f[284] && !f[145];
	assign leaf[1216] = f[154] && f[577] && !f[284] && f[145];
	assign leaf[1217] = f[154] && f[577] && f[284];
	
	// Tree 78, Classifier 8, Iteration: 7
	assign leaf[1218] = !f[658] && !f[652] && !f[686] && !f[303];
	assign leaf[1219] = !f[658] && !f[652] && !f[686] && f[303];
	assign leaf[1220] = !f[658] && !f[652] && f[686] && !f[571];
	assign leaf[1221] = !f[658] && !f[652] && f[686] && f[571];
	assign leaf[1222] = !f[658] && f[652] && !f[513] && !f[599];
	assign leaf[1223] = !f[658] && f[652] && !f[513] && f[599];
	assign leaf[1224] = !f[658] && f[652] && f[513] && !f[570];
	assign leaf[1225] = !f[658] && f[652] && f[513] && f[570];
	assign leaf[1226] = f[658] && !f[543] && !f[541] && !f[544];
	assign leaf[1227] = f[658] && !f[543] && !f[541] && f[544];
	assign leaf[1228] = f[658] && !f[543] && f[541] && !f[379];
	assign leaf[1229] = f[658] && !f[543] && f[541] && f[379];
	assign leaf[1230] = f[658] && f[543] && !f[484] && !f[601];
	assign leaf[1231] = f[658] && f[543] && !f[484] && f[601];
	assign leaf[1232] = f[658] && f[543] && f[484] && !f[303];
	assign leaf[1233] = f[658] && f[543] && f[484] && f[303];
	
	// Tree 79, Classifier 9, Iteration: 7
	assign leaf[1234] = !f[570] && !f[624] && !f[212] && !f[719];
	assign leaf[1235] = !f[570] && !f[624] && !f[212] && f[719];
	assign leaf[1236] = !f[570] && !f[624] && f[212] && !f[204];
	assign leaf[1237] = !f[570] && !f[624] && f[212] && f[204];
	assign leaf[1238] = !f[570] && f[624] && !f[384] && !f[324];
	assign leaf[1239] = !f[570] && f[624] && !f[384] && f[324];
	assign leaf[1240] = !f[570] && f[624] && f[384] && !f[680];
	assign leaf[1241] = !f[570] && f[624] && f[384] && f[680];
	assign leaf[1242] = f[570] && !f[680] && !f[720] && !f[599];
	assign leaf[1243] = f[570] && !f[680] && !f[720] && f[599];
	assign leaf[1244] = f[570] && !f[680] && f[720];
	assign leaf[1245] = f[570] && f[680] && !f[207] && !f[213];
	assign leaf[1246] = f[570] && f[680] && !f[207] && f[213];
	assign leaf[1247] = f[570] && f[680] && f[207] && !f[377];
	assign leaf[1248] = f[570] && f[680] && f[207] && f[377];
	
	// Tree 80, Classifier 0, Iteration: 8
	assign leaf[1249] = !f[408] && !f[427] && !f[429] && !f[425];
	assign leaf[1250] = !f[408] && !f[427] && !f[429] && f[425];
	assign leaf[1251] = !f[408] && !f[427] && f[429] && !f[485];
	assign leaf[1252] = !f[408] && !f[427] && f[429] && f[485];
	assign leaf[1253] = !f[408] && f[427] && !f[460] && !f[716];
	assign leaf[1254] = !f[408] && f[427] && !f[460] && f[716];
	assign leaf[1255] = !f[408] && f[427] && f[460] && !f[292];
	assign leaf[1256] = !f[408] && f[427] && f[460] && f[292];
	assign leaf[1257] = f[408] && !f[293] && !f[455];
	assign leaf[1258] = f[408] && !f[293] && f[455] && !f[656];
	assign leaf[1259] = f[408] && !f[293] && f[455] && f[656];
	assign leaf[1260] = f[408] && f[293] && !f[406] && !f[404];
	assign leaf[1261] = f[408] && f[293] && !f[406] && f[404];
	assign leaf[1262] = f[408] && f[293] && f[406] && !f[414];
	assign leaf[1263] = f[408] && f[293] && f[406] && f[414];
	
	// Tree 81, Classifier 1, Iteration: 8
	assign leaf[1264] = !f[402] && !f[406] && !f[99] && !f[405];
	assign leaf[1265] = !f[402] && !f[406] && !f[99] && f[405];
	assign leaf[1266] = !f[402] && !f[406] && f[99] && !f[379];
	assign leaf[1267] = !f[402] && !f[406] && f[99] && f[379];
	assign leaf[1268] = !f[402] && f[406] && !f[233] && !f[295];
	assign leaf[1269] = !f[402] && f[406] && !f[233] && f[295];
	assign leaf[1270] = !f[402] && f[406] && f[233] && !f[269];
	assign leaf[1271] = !f[402] && f[406] && f[233] && f[269];
	assign leaf[1272] = f[402] && !f[295];
	assign leaf[1273] = f[402] && f[295] && !f[494] && !f[373];
	assign leaf[1274] = f[402] && f[295] && !f[494] && f[373];
	assign leaf[1275] = f[402] && f[295] && f[494];
	
	// Tree 82, Classifier 2, Iteration: 8
	assign leaf[1276] = !f[543] && !f[125] && !f[511] && !f[501];
	assign leaf[1277] = !f[543] && !f[125] && !f[511] && f[501];
	assign leaf[1278] = !f[543] && !f[125] && f[511] && !f[630];
	assign leaf[1279] = !f[543] && !f[125] && f[511] && f[630];
	assign leaf[1280] = !f[543] && f[125] && !f[458] && !f[631];
	assign leaf[1281] = !f[543] && f[125] && !f[458] && f[631];
	assign leaf[1282] = !f[543] && f[125] && f[458] && !f[659];
	assign leaf[1283] = !f[543] && f[125] && f[458] && f[659];
	assign leaf[1284] = f[543] && !f[607] && !f[524] && !f[470];
	assign leaf[1285] = f[543] && !f[607] && !f[524] && f[470];
	assign leaf[1286] = f[543] && !f[607] && f[524] && !f[344];
	assign leaf[1287] = f[543] && !f[607] && f[524] && f[344];
	assign leaf[1288] = f[543] && f[607] && !f[496] && !f[442];
	assign leaf[1289] = f[543] && f[607] && !f[496] && f[442];
	assign leaf[1290] = f[543] && f[607] && f[496] && !f[594];
	assign leaf[1291] = f[543] && f[607] && f[496] && f[594];
	
	// Tree 83, Classifier 3, Iteration: 8
	assign leaf[1292] = !f[655] && !f[710] && !f[627] && !f[175];
	assign leaf[1293] = !f[655] && !f[710] && !f[627] && f[175];
	assign leaf[1294] = !f[655] && !f[710] && f[627] && !f[457];
	assign leaf[1295] = !f[655] && !f[710] && f[627] && f[457];
	assign leaf[1296] = !f[655] && f[710] && !f[485] && !f[265];
	assign leaf[1297] = !f[655] && f[710] && !f[485] && f[265];
	assign leaf[1298] = !f[655] && f[710] && f[485];
	assign leaf[1299] = f[655] && !f[517] && !f[318] && !f[343];
	assign leaf[1300] = f[655] && !f[517] && !f[318] && f[343];
	assign leaf[1301] = f[655] && !f[517] && f[318] && !f[148];
	assign leaf[1302] = f[655] && !f[517] && f[318] && f[148];
	assign leaf[1303] = f[655] && f[517] && !f[603] && !f[153];
	assign leaf[1304] = f[655] && f[517] && !f[603] && f[153];
	assign leaf[1305] = f[655] && f[517] && f[603] && !f[290];
	assign leaf[1306] = f[655] && f[517] && f[603] && f[290];
	
	// Tree 84, Classifier 4, Iteration: 8
	assign leaf[1307] = !f[568] && !f[455] && !f[238] && !f[182];
	assign leaf[1308] = !f[568] && !f[455] && !f[238] && f[182];
	assign leaf[1309] = !f[568] && !f[455] && f[238] && !f[240];
	assign leaf[1310] = !f[568] && !f[455] && f[238] && f[240];
	assign leaf[1311] = !f[568] && f[455] && !f[347] && !f[238];
	assign leaf[1312] = !f[568] && f[455] && !f[347] && f[238];
	assign leaf[1313] = !f[568] && f[455] && f[347] && !f[491];
	assign leaf[1314] = !f[568] && f[455] && f[347] && f[491];
	assign leaf[1315] = f[568] && !f[626] && !f[135] && !f[381];
	assign leaf[1316] = f[568] && !f[626] && !f[135] && f[381];
	assign leaf[1317] = f[568] && !f[626] && f[135] && !f[598];
	assign leaf[1318] = f[568] && !f[626] && f[135] && f[598];
	assign leaf[1319] = f[568] && f[626] && !f[426] && !f[136];
	assign leaf[1320] = f[568] && f[626] && !f[426] && f[136];
	assign leaf[1321] = f[568] && f[626] && f[426] && !f[462];
	assign leaf[1322] = f[568] && f[626] && f[426] && f[462];
	
	// Tree 85, Classifier 5, Iteration: 8
	assign leaf[1323] = !f[488] && !f[188] && !f[247] && !f[158];
	assign leaf[1324] = !f[488] && !f[188] && !f[247] && f[158];
	assign leaf[1325] = !f[488] && !f[188] && f[247] && !f[356];
	assign leaf[1326] = !f[488] && !f[188] && f[247] && f[356];
	assign leaf[1327] = !f[488] && f[188] && !f[272] && !f[303];
	assign leaf[1328] = !f[488] && f[188] && !f[272] && f[303];
	assign leaf[1329] = !f[488] && f[188] && f[272] && !f[219];
	assign leaf[1330] = !f[488] && f[188] && f[272] && f[219];
	assign leaf[1331] = f[488] && !f[380] && !f[410] && !f[374];
	assign leaf[1332] = f[488] && !f[380] && !f[410] && f[374];
	assign leaf[1333] = f[488] && !f[380] && f[410] && !f[583];
	assign leaf[1334] = f[488] && !f[380] && f[410] && f[583];
	assign leaf[1335] = f[488] && f[380] && !f[461] && !f[245];
	assign leaf[1336] = f[488] && f[380] && !f[461] && f[245];
	assign leaf[1337] = f[488] && f[380] && f[461] && !f[353];
	assign leaf[1338] = f[488] && f[380] && f[461] && f[353];
	
	// Tree 86, Classifier 6, Iteration: 8
	assign leaf[1339] = !f[486] && !f[484] && !f[388] && !f[487];
	assign leaf[1340] = !f[486] && !f[484] && !f[388] && f[487];
	assign leaf[1341] = !f[486] && !f[484] && f[388] && !f[266];
	assign leaf[1342] = !f[486] && !f[484] && f[388] && f[266];
	assign leaf[1343] = !f[486] && f[484] && !f[243] && !f[217];
	assign leaf[1344] = !f[486] && f[484] && !f[243] && f[217];
	assign leaf[1345] = !f[486] && f[484] && f[243] && !f[93];
	assign leaf[1346] = !f[486] && f[484] && f[243] && f[93];
	assign leaf[1347] = f[486] && !f[271] && !f[402] && !f[414];
	assign leaf[1348] = f[486] && !f[271] && !f[402] && f[414];
	assign leaf[1349] = f[486] && !f[271] && f[402] && !f[274];
	assign leaf[1350] = f[486] && !f[271] && f[402] && f[274];
	assign leaf[1351] = f[486] && f[271] && !f[121] && !f[96];
	assign leaf[1352] = f[486] && f[271] && !f[121] && f[96];
	assign leaf[1353] = f[486] && f[271] && f[121] && !f[185];
	assign leaf[1354] = f[486] && f[271] && f[121] && f[185];
	
	// Tree 87, Classifier 7, Iteration: 8
	assign leaf[1355] = !f[267] && !f[745] && !f[402] && !f[377];
	assign leaf[1356] = !f[267] && !f[745] && !f[402] && f[377];
	assign leaf[1357] = !f[267] && !f[745] && f[402] && !f[295];
	assign leaf[1358] = !f[267] && !f[745] && f[402] && f[295];
	assign leaf[1359] = !f[267] && f[745] && !f[432] && !f[373];
	assign leaf[1360] = !f[267] && f[745] && !f[432] && f[373];
	assign leaf[1361] = !f[267] && f[745] && f[432];
	assign leaf[1362] = f[267] && !f[263] && !f[236] && !f[290];
	assign leaf[1363] = f[267] && !f[263] && !f[236] && f[290];
	assign leaf[1364] = f[267] && !f[263] && f[236] && !f[606];
	assign leaf[1365] = f[267] && !f[263] && f[236] && f[606];
	assign leaf[1366] = f[267] && f[263] && !f[567] && !f[403];
	assign leaf[1367] = f[267] && f[263] && !f[567] && f[403];
	assign leaf[1368] = f[267] && f[263] && f[567] && !f[677];
	assign leaf[1369] = f[267] && f[263] && f[567] && f[677];
	
	// Tree 88, Classifier 8, Iteration: 8
	assign leaf[1370] = !f[439] && !f[267] && !f[349] && !f[375];
	assign leaf[1371] = !f[439] && !f[267] && !f[349] && f[375];
	assign leaf[1372] = !f[439] && !f[267] && f[349] && !f[406];
	assign leaf[1373] = !f[439] && !f[267] && f[349] && f[406];
	assign leaf[1374] = !f[439] && f[267] && !f[301] && !f[661];
	assign leaf[1375] = !f[439] && f[267] && !f[301] && f[661];
	assign leaf[1376] = !f[439] && f[267] && f[301] && !f[380];
	assign leaf[1377] = !f[439] && f[267] && f[301] && f[380];
	assign leaf[1378] = f[439] && !f[521] && !f[330] && !f[377];
	assign leaf[1379] = f[439] && !f[521] && !f[330] && f[377];
	assign leaf[1380] = f[439] && !f[521] && f[330] && !f[355];
	assign leaf[1381] = f[439] && !f[521] && f[330] && f[355];
	assign leaf[1382] = f[439] && f[521] && !f[304] && !f[154];
	assign leaf[1383] = f[439] && f[521] && !f[304] && f[154];
	assign leaf[1384] = f[439] && f[521] && f[304] && !f[468];
	assign leaf[1385] = f[439] && f[521] && f[304] && f[468];
	
	// Tree 89, Classifier 9, Iteration: 8
	assign leaf[1386] = !f[157] && !f[571] && !f[203] && !f[189];
	assign leaf[1387] = !f[157] && !f[571] && !f[203] && f[189];
	assign leaf[1388] = !f[157] && !f[571] && f[203] && !f[342];
	assign leaf[1389] = !f[157] && !f[571] && f[203] && f[342];
	assign leaf[1390] = !f[157] && f[571] && !f[709] && !f[679];
	assign leaf[1391] = !f[157] && f[571] && !f[709] && f[679];
	assign leaf[1392] = !f[157] && f[571] && f[709] && !f[185];
	assign leaf[1393] = !f[157] && f[571] && f[709] && f[185];
	assign leaf[1394] = f[157] && !f[372] && !f[397] && !f[291];
	assign leaf[1395] = f[157] && !f[372] && !f[397] && f[291];
	assign leaf[1396] = f[157] && !f[372] && f[397] && !f[552];
	assign leaf[1397] = f[157] && !f[372] && f[397] && f[552];
	assign leaf[1398] = f[157] && f[372] && !f[235] && !f[236];
	assign leaf[1399] = f[157] && f[372] && !f[235] && f[236];
	assign leaf[1400] = f[157] && f[372] && f[235] && !f[552];
	assign leaf[1401] = f[157] && f[372] && f[235] && f[552];
	
	// Tree 90, Classifier 0, Iteration: 9
	assign leaf[1402] = !f[462] && !f[378] && !f[402] && !f[410];
	assign leaf[1403] = !f[462] && !f[378] && !f[402] && f[410];
	assign leaf[1404] = !f[462] && !f[378] && f[402] && !f[599];
	assign leaf[1405] = !f[462] && !f[378] && f[402] && f[599];
	assign leaf[1406] = !f[462] && f[378] && !f[273] && !f[274];
	assign leaf[1407] = !f[462] && f[378] && !f[273] && f[274];
	assign leaf[1408] = !f[462] && f[378] && f[273] && !f[266];
	assign leaf[1409] = !f[462] && f[378] && f[273] && f[266];
	assign leaf[1410] = f[462] && !f[386] && !f[568] && !f[508];
	assign leaf[1411] = f[462] && !f[386] && !f[568] && f[508];
	assign leaf[1412] = f[462] && !f[386] && f[568] && !f[461];
	assign leaf[1413] = f[462] && !f[386] && f[568] && f[461];
	assign leaf[1414] = f[462] && f[386] && !f[297] && !f[273];
	assign leaf[1415] = f[462] && f[386] && !f[297] && f[273];
	assign leaf[1416] = f[462] && f[386] && f[297] && !f[155];
	assign leaf[1417] = f[462] && f[386] && f[297] && f[155];
	
	// Tree 91, Classifier 1, Iteration: 9
	assign leaf[1418] = !f[410] && !f[318] && !f[511] && !f[205];
	assign leaf[1419] = !f[410] && !f[318] && !f[511] && f[205];
	assign leaf[1420] = !f[410] && !f[318] && f[511] && !f[649];
	assign leaf[1421] = !f[410] && !f[318] && f[511] && f[649];
	assign leaf[1422] = !f[410] && f[318] && !f[294] && !f[148];
	assign leaf[1423] = !f[410] && f[318] && !f[294] && f[148];
	assign leaf[1424] = !f[410] && f[318] && f[294] && !f[126];
	assign leaf[1425] = !f[410] && f[318] && f[294] && f[126];
	assign leaf[1426] = f[410] && !f[163] && !f[411] && !f[322];
	assign leaf[1427] = f[410] && !f[163] && !f[411] && f[322];
	assign leaf[1428] = f[410] && !f[163] && f[411];
	assign leaf[1429] = f[410] && f[163] && !f[269];
	assign leaf[1430] = f[410] && f[163] && f[269];
	
	// Tree 92, Classifier 2, Iteration: 9
	assign leaf[1431] = !f[345] && !f[320] && !f[343] && !f[379];
	assign leaf[1432] = !f[345] && !f[320] && !f[343] && f[379];
	assign leaf[1433] = !f[345] && !f[320] && f[343] && !f[399];
	assign leaf[1434] = !f[345] && !f[320] && f[343] && f[399];
	assign leaf[1435] = !f[345] && f[320] && !f[554] && !f[473];
	assign leaf[1436] = !f[345] && f[320] && !f[554] && f[473];
	assign leaf[1437] = !f[345] && f[320] && f[554] && !f[660];
	assign leaf[1438] = !f[345] && f[320] && f[554] && f[660];
	assign leaf[1439] = f[345] && !f[568] && !f[401] && !f[515];
	assign leaf[1440] = f[345] && !f[568] && !f[401] && f[515];
	assign leaf[1441] = f[345] && !f[568] && f[401] && !f[511];
	assign leaf[1442] = f[345] && !f[568] && f[401] && f[511];
	assign leaf[1443] = f[345] && f[568] && !f[464] && !f[622];
	assign leaf[1444] = f[345] && f[568] && !f[464] && f[622];
	assign leaf[1445] = f[345] && f[568] && f[464] && !f[658];
	assign leaf[1446] = f[345] && f[568] && f[464] && f[658];
	
	// Tree 93, Classifier 3, Iteration: 9
	assign leaf[1447] = !f[518] && !f[344] && !f[516] && !f[485];
	assign leaf[1448] = !f[518] && !f[344] && !f[516] && f[485];
	assign leaf[1449] = !f[518] && !f[344] && f[516] && !f[488];
	assign leaf[1450] = !f[518] && !f[344] && f[516] && f[488];
	assign leaf[1451] = !f[518] && f[344] && !f[288] && !f[348];
	assign leaf[1452] = !f[518] && f[344] && !f[288] && f[348];
	assign leaf[1453] = !f[518] && f[344] && f[288] && !f[291];
	assign leaf[1454] = !f[518] && f[344] && f[288] && f[291];
	assign leaf[1455] = f[518] && !f[463] && !f[352] && !f[632];
	assign leaf[1456] = f[518] && !f[463] && !f[352] && f[632];
	assign leaf[1457] = f[518] && !f[463] && f[352] && !f[373];
	assign leaf[1458] = f[518] && !f[463] && f[352] && f[373];
	assign leaf[1459] = f[518] && f[463] && !f[623] && !f[536];
	assign leaf[1460] = f[518] && f[463] && !f[623] && f[536];
	assign leaf[1461] = f[518] && f[463] && f[623] && !f[352];
	assign leaf[1462] = f[518] && f[463] && f[623] && f[352];
	
	// Tree 94, Classifier 4, Iteration: 9
	assign leaf[1463] = !f[464] && !f[603] && !f[295] && !f[659];
	assign leaf[1464] = !f[464] && !f[603] && !f[295] && f[659];
	assign leaf[1465] = !f[464] && !f[603] && f[295] && !f[346];
	assign leaf[1466] = !f[464] && !f[603] && f[295] && f[346];
	assign leaf[1467] = !f[464] && f[603] && !f[688] && !f[686];
	assign leaf[1468] = !f[464] && f[603] && !f[688] && f[686];
	assign leaf[1469] = !f[464] && f[603] && f[688] && !f[210];
	assign leaf[1470] = !f[464] && f[603] && f[688] && f[210];
	assign leaf[1471] = f[464] && !f[569] && !f[208] && !f[710];
	assign leaf[1472] = f[464] && !f[569] && !f[208] && f[710];
	assign leaf[1473] = f[464] && !f[569] && f[208] && !f[319];
	assign leaf[1474] = f[464] && !f[569] && f[208] && f[319];
	assign leaf[1475] = f[464] && f[569] && !f[163] && !f[399];
	assign leaf[1476] = f[464] && f[569] && !f[163] && f[399];
	assign leaf[1477] = f[464] && f[569] && f[163] && !f[213];
	assign leaf[1478] = f[464] && f[569] && f[163] && f[213];
	
	// Tree 95, Classifier 5, Iteration: 9
	assign leaf[1479] = !f[463] && !f[269] && !f[266] && !f[271];
	assign leaf[1480] = !f[463] && !f[269] && !f[266] && f[271];
	assign leaf[1481] = !f[463] && !f[269] && f[266] && !f[215];
	assign leaf[1482] = !f[463] && !f[269] && f[266] && f[215];
	assign leaf[1483] = !f[463] && f[269] && !f[245] && !f[305];
	assign leaf[1484] = !f[463] && f[269] && !f[245] && f[305];
	assign leaf[1485] = !f[463] && f[269] && f[245] && !f[386];
	assign leaf[1486] = !f[463] && f[269] && f[245] && f[386];
	assign leaf[1487] = f[463] && !f[353] && !f[383] && !f[351];
	assign leaf[1488] = f[463] && !f[353] && !f[383] && f[351];
	assign leaf[1489] = f[463] && !f[353] && f[383] && !f[525];
	assign leaf[1490] = f[463] && !f[353] && f[383] && f[525];
	assign leaf[1491] = f[463] && f[353] && !f[304] && !f[322];
	assign leaf[1492] = f[463] && f[353] && !f[304] && f[322];
	assign leaf[1493] = f[463] && f[353] && f[304] && !f[213];
	assign leaf[1494] = f[463] && f[353] && f[304] && f[213];
	
	// Tree 96, Classifier 6, Iteration: 9
	assign leaf[1495] = !f[269] && !f[244] && !f[323] && !f[246];
	assign leaf[1496] = !f[269] && !f[244] && !f[323] && f[246];
	assign leaf[1497] = !f[269] && !f[244] && f[323] && !f[430];
	assign leaf[1498] = !f[269] && !f[244] && f[323] && f[430];
	assign leaf[1499] = !f[269] && f[244] && !f[355] && !f[513];
	assign leaf[1500] = !f[269] && f[244] && !f[355] && f[513];
	assign leaf[1501] = !f[269] && f[244] && f[355] && !f[414];
	assign leaf[1502] = !f[269] && f[244] && f[355] && f[414];
	assign leaf[1503] = f[269] && !f[133] && !f[386] && !f[164];
	assign leaf[1504] = f[269] && !f[133] && !f[386] && f[164];
	assign leaf[1505] = f[269] && !f[133] && f[386] && !f[239];
	assign leaf[1506] = f[269] && !f[133] && f[386] && f[239];
	assign leaf[1507] = f[269] && f[133] && !f[325] && !f[273];
	assign leaf[1508] = f[269] && f[133] && !f[325] && f[273];
	assign leaf[1509] = f[269] && f[133] && f[325] && !f[266];
	assign leaf[1510] = f[269] && f[133] && f[325] && f[266];
	
	// Tree 97, Classifier 7, Iteration: 9
	assign leaf[1511] = !f[157] && !f[376] && !f[552] && !f[401];
	assign leaf[1512] = !f[157] && !f[376] && !f[552] && f[401];
	assign leaf[1513] = !f[157] && !f[376] && f[552] && !f[746];
	assign leaf[1514] = !f[157] && !f[376] && f[552] && f[746];
	assign leaf[1515] = !f[157] && f[376] && !f[340] && !f[411];
	assign leaf[1516] = !f[157] && f[376] && !f[340] && f[411];
	assign leaf[1517] = !f[157] && f[376] && f[340] && !f[430];
	assign leaf[1518] = !f[157] && f[376] && f[340] && f[430];
	assign leaf[1519] = f[157] && !f[518];
	assign leaf[1520] = f[157] && f[518] && !f[148] && !f[685];
	assign leaf[1521] = f[157] && f[518] && !f[148] && f[685];
	assign leaf[1522] = f[157] && f[518] && f[148] && !f[552];
	assign leaf[1523] = f[157] && f[518] && f[148] && f[552];
	
	// Tree 98, Classifier 8, Iteration: 9
	assign leaf[1524] = !f[658] && !f[624] && !f[686] && !f[630];
	assign leaf[1525] = !f[658] && !f[624] && !f[686] && f[630];
	assign leaf[1526] = !f[658] && !f[624] && f[686] && !f[516];
	assign leaf[1527] = !f[658] && !f[624] && f[686] && f[516];
	assign leaf[1528] = !f[658] && f[624] && !f[571] && !f[494];
	assign leaf[1529] = !f[658] && f[624] && !f[571] && f[494];
	assign leaf[1530] = !f[658] && f[624] && f[571] && !f[265];
	assign leaf[1531] = !f[658] && f[624] && f[571] && f[265];
	assign leaf[1532] = f[658] && !f[516] && !f[513] && !f[511];
	assign leaf[1533] = f[658] && !f[516] && !f[513] && f[511];
	assign leaf[1534] = f[658] && !f[516] && f[513] && !f[379];
	assign leaf[1535] = f[658] && !f[516] && f[513] && f[379];
	assign leaf[1536] = f[658] && f[516] && !f[602] && !f[514];
	assign leaf[1537] = f[658] && f[516] && !f[602] && f[514];
	assign leaf[1538] = f[658] && f[516] && f[602] && !f[317];
	assign leaf[1539] = f[658] && f[516] && f[602] && f[317];
	
	// Tree 99, Classifier 9, Iteration: 9
	assign leaf[1540] = !f[154] && !f[596] && !f[210] && !f[266];
	assign leaf[1541] = !f[154] && !f[596] && !f[210] && f[266];
	assign leaf[1542] = !f[154] && !f[596] && f[210] && !f[206];
	assign leaf[1543] = !f[154] && !f[596] && f[210] && f[206];
	assign leaf[1544] = !f[154] && f[596] && !f[706] && !f[665];
	assign leaf[1545] = !f[154] && f[596] && !f[706] && f[665];
	assign leaf[1546] = !f[154] && f[596] && f[706] && !f[375];
	assign leaf[1547] = !f[154] && f[596] && f[706] && f[375];
	assign leaf[1548] = f[154] && !f[316] && !f[290] && !f[342];
	assign leaf[1549] = f[154] && !f[316] && !f[290] && f[342];
	assign leaf[1550] = f[154] && !f[316] && f[290] && !f[571];
	assign leaf[1551] = f[154] && !f[316] && f[290] && f[571];
	assign leaf[1552] = f[154] && f[316] && !f[600] && !f[354];
	assign leaf[1553] = f[154] && f[316] && !f[600] && f[354];
	assign leaf[1554] = f[154] && f[316] && f[600] && !f[544];
	assign leaf[1555] = f[154] && f[316] && f[600] && f[544];
	
	// Tree 100, Classifier 0, Iteration: 10
	assign leaf[1556] = !f[434] && !f[455] && !f[458] && !f[425];
	assign leaf[1557] = !f[434] && !f[455] && !f[458] && f[425];
	assign leaf[1558] = !f[434] && !f[455] && f[458] && !f[355];
	assign leaf[1559] = !f[434] && !f[455] && f[458] && f[355];
	assign leaf[1560] = !f[434] && f[455] && !f[539] && !f[437];
	assign leaf[1561] = !f[434] && f[455] && !f[539] && f[437];
	assign leaf[1562] = !f[434] && f[455] && f[539] && !f[98];
	assign leaf[1563] = !f[434] && f[455] && f[539] && f[98];
	assign leaf[1564] = f[434] && !f[385] && !f[360] && !f[383];
	assign leaf[1565] = f[434] && !f[385] && !f[360] && f[383];
	assign leaf[1566] = f[434] && !f[385] && f[360];
	assign leaf[1567] = f[434] && f[385] && !f[468] && !f[536];
	assign leaf[1568] = f[434] && f[385] && !f[468] && f[536];
	assign leaf[1569] = f[434] && f[385] && f[468] && !f[213];
	assign leaf[1570] = f[434] && f[385] && f[468] && f[213];
	
	// Tree 101, Classifier 1, Iteration: 10
	assign leaf[1571] = !f[430] && !f[434] && !f[433] && !f[101];
	assign leaf[1572] = !f[430] && !f[434] && !f[433] && f[101];
	assign leaf[1573] = !f[430] && !f[434] && f[433] && !f[548];
	assign leaf[1574] = !f[430] && !f[434] && f[433] && f[548];
	assign leaf[1575] = !f[430] && f[434] && !f[299] && !f[322];
	assign leaf[1576] = !f[430] && f[434] && !f[299] && f[322];
	assign leaf[1577] = !f[430] && f[434] && f[299] && !f[183];
	assign leaf[1578] = !f[430] && f[434] && f[299] && f[183];
	assign leaf[1579] = f[430] && !f[349] && !f[649] && !f[743];
	assign leaf[1580] = f[430] && !f[349] && !f[649] && f[743];
	assign leaf[1581] = f[430] && !f[349] && f[649] && !f[184];
	assign leaf[1582] = f[430] && !f[349] && f[649] && f[184];
	assign leaf[1583] = f[430] && f[349] && !f[521] && !f[268];
	assign leaf[1584] = f[430] && f[349] && !f[521] && f[268];
	assign leaf[1585] = f[430] && f[349] && f[521];
	
	// Tree 102, Classifier 2, Iteration: 10
	assign leaf[1586] = !f[151] && !f[657] && !f[156] && !f[527];
	assign leaf[1587] = !f[151] && !f[657] && !f[156] && f[527];
	assign leaf[1588] = !f[151] && !f[657] && f[156] && !f[322];
	assign leaf[1589] = !f[151] && !f[657] && f[156] && f[322];
	assign leaf[1590] = !f[151] && f[657] && !f[636] && !f[717];
	assign leaf[1591] = !f[151] && f[657] && !f[636] && f[717];
	assign leaf[1592] = !f[151] && f[657] && f[636] && !f[516];
	assign leaf[1593] = !f[151] && f[657] && f[636] && f[516];
	assign leaf[1594] = f[151] && !f[317] && !f[545] && !f[487];
	assign leaf[1595] = f[151] && !f[317] && !f[545] && f[487];
	assign leaf[1596] = f[151] && !f[317] && f[545] && !f[342];
	assign leaf[1597] = f[151] && !f[317] && f[545] && f[342];
	assign leaf[1598] = f[151] && f[317] && !f[639] && !f[372];
	assign leaf[1599] = f[151] && f[317] && !f[639] && f[372];
	assign leaf[1600] = f[151] && f[317] && f[639] && !f[554];
	assign leaf[1601] = f[151] && f[317] && f[639] && f[554];
	
	// Tree 103, Classifier 3, Iteration: 10
	assign leaf[1602] = !f[655] && !f[400] && !f[495] && !f[469];
	assign leaf[1603] = !f[655] && !f[400] && !f[495] && f[469];
	assign leaf[1604] = !f[655] && !f[400] && f[495] && !f[458];
	assign leaf[1605] = !f[655] && !f[400] && f[495] && f[458];
	assign leaf[1606] = !f[655] && f[400] && !f[200] && !f[710];
	assign leaf[1607] = !f[655] && f[400] && !f[200] && f[710];
	assign leaf[1608] = !f[655] && f[400] && f[200] && !f[314];
	assign leaf[1609] = !f[655] && f[400] && f[200] && f[314];
	assign leaf[1610] = f[655] && !f[291] && !f[544] && !f[317];
	assign leaf[1611] = f[655] && !f[291] && !f[544] && f[317];
	assign leaf[1612] = f[655] && !f[291] && f[544] && !f[489];
	assign leaf[1613] = f[655] && !f[291] && f[544] && f[489];
	assign leaf[1614] = f[655] && f[291] && !f[149] && !f[319];
	assign leaf[1615] = f[655] && f[291] && !f[149] && f[319];
	assign leaf[1616] = f[655] && f[291] && f[149] && !f[261];
	assign leaf[1617] = f[655] && f[291] && f[149] && f[261];
	
	// Tree 104, Classifier 4, Iteration: 10
	assign leaf[1618] = !f[463] && !f[628] && !f[322] && !f[238];
	assign leaf[1619] = !f[463] && !f[628] && !f[322] && f[238];
	assign leaf[1620] = !f[463] && !f[628] && f[322] && !f[375];
	assign leaf[1621] = !f[463] && !f[628] && f[322] && f[375];
	assign leaf[1622] = !f[463] && f[628] && !f[163] && !f[490];
	assign leaf[1623] = !f[463] && f[628] && !f[163] && f[490];
	assign leaf[1624] = !f[463] && f[628] && f[163] && !f[595];
	assign leaf[1625] = !f[463] && f[628] && f[163] && f[595];
	assign leaf[1626] = f[463] && !f[542] && !f[624] && !f[347];
	assign leaf[1627] = f[463] && !f[542] && !f[624] && f[347];
	assign leaf[1628] = f[463] && !f[542] && f[624] && !f[516];
	assign leaf[1629] = f[463] && !f[542] && f[624] && f[516];
	assign leaf[1630] = f[463] && f[542] && !f[163] && !f[220];
	assign leaf[1631] = f[463] && f[542] && !f[163] && f[220];
	assign leaf[1632] = f[463] && f[542] && f[163] && !f[213];
	assign leaf[1633] = f[463] && f[542] && f[163] && f[213];
	
	// Tree 105, Classifier 5, Iteration: 10
	assign leaf[1634] = !f[487] && !f[598] && !f[546] && !f[296];
	assign leaf[1635] = !f[487] && !f[598] && !f[546] && f[296];
	assign leaf[1636] = !f[487] && !f[598] && f[546] && !f[542];
	assign leaf[1637] = !f[487] && !f[598] && f[546] && f[542];
	assign leaf[1638] = !f[487] && f[598] && !f[456] && !f[133];
	assign leaf[1639] = !f[487] && f[598] && !f[456] && f[133];
	assign leaf[1640] = !f[487] && f[598] && f[456] && !f[484];
	assign leaf[1641] = !f[487] && f[598] && f[456] && f[484];
	assign leaf[1642] = f[487] && !f[247] && !f[660] && !f[275];
	assign leaf[1643] = f[487] && !f[247] && !f[660] && f[275];
	assign leaf[1644] = f[487] && !f[247] && f[660] && !f[297];
	assign leaf[1645] = f[487] && !f[247] && f[660] && f[297];
	assign leaf[1646] = f[487] && f[247] && !f[356] && !f[268];
	assign leaf[1647] = f[487] && f[247] && !f[356] && f[268];
	assign leaf[1648] = f[487] && f[247] && f[356] && !f[710];
	assign leaf[1649] = f[487] && f[247] && f[356] && f[710];
	
	// Tree 106, Classifier 6, Iteration: 10
	assign leaf[1650] = !f[269] && !f[243] && !f[549] && !f[323];
	assign leaf[1651] = !f[269] && !f[243] && !f[549] && f[323];
	assign leaf[1652] = !f[269] && !f[243] && f[549] && !f[633];
	assign leaf[1653] = !f[269] && !f[243] && f[549] && f[633];
	assign leaf[1654] = !f[269] && f[243] && !f[327] && !f[486];
	assign leaf[1655] = !f[269] && f[243] && !f[327] && f[486];
	assign leaf[1656] = !f[269] && f[243] && f[327] && !f[358];
	assign leaf[1657] = !f[269] && f[243] && f[327] && f[358];
	assign leaf[1658] = f[269] && !f[133] && !f[94] && !f[103];
	assign leaf[1659] = f[269] && !f[133] && !f[94] && f[103];
	assign leaf[1660] = f[269] && !f[133] && f[94] && !f[232];
	assign leaf[1661] = f[269] && !f[133] && f[94] && f[232];
	assign leaf[1662] = f[269] && f[133] && !f[299] && !f[349];
	assign leaf[1663] = f[269] && f[133] && !f[299] && f[349];
	assign leaf[1664] = f[269] && f[133] && f[299];
	
	// Tree 107, Classifier 7, Iteration: 10
	assign leaf[1665] = !f[154] && !f[159] && !f[432] && !f[486];
	assign leaf[1666] = !f[154] && !f[159] && !f[432] && f[486];
	assign leaf[1667] = !f[154] && !f[159] && f[432] && !f[345];
	assign leaf[1668] = !f[154] && !f[159] && f[432] && f[345];
	assign leaf[1669] = !f[154] && f[159] && !f[206];
	assign leaf[1670] = !f[154] && f[159] && f[206] && !f[268];
	assign leaf[1671] = !f[154] && f[159] && f[206] && f[268];
	assign leaf[1672] = f[154] && !f[577] && !f[679] && !f[240];
	assign leaf[1673] = f[154] && !f[577] && !f[679] && f[240];
	assign leaf[1674] = f[154] && !f[577] && f[679] && !f[377];
	assign leaf[1675] = f[154] && !f[577] && f[679] && f[377];
	assign leaf[1676] = f[154] && f[577] && !f[145];
	assign leaf[1677] = f[154] && f[577] && f[145];
	
	// Tree 108, Classifier 8, Iteration: 10
	assign leaf[1678] = !f[439] && !f[302] && !f[183] && !f[154];
	assign leaf[1679] = !f[439] && !f[302] && !f[183] && f[154];
	assign leaf[1680] = !f[439] && !f[302] && f[183] && !f[299];
	assign leaf[1681] = !f[439] && !f[302] && f[183] && f[299];
	assign leaf[1682] = !f[439] && f[302] && !f[469] && !f[272];
	assign leaf[1683] = !f[439] && f[302] && !f[469] && f[272];
	assign leaf[1684] = !f[439] && f[302] && f[469] && !f[399];
	assign leaf[1685] = !f[439] && f[302] && f[469] && f[399];
	assign leaf[1686] = f[439] && !f[521] && !f[179] && !f[331];
	assign leaf[1687] = f[439] && !f[521] && !f[179] && f[331];
	assign leaf[1688] = f[439] && !f[521] && f[179] && !f[550];
	assign leaf[1689] = f[439] && !f[521] && f[179] && f[550];
	assign leaf[1690] = f[439] && f[521] && !f[304] && !f[378];
	assign leaf[1691] = f[439] && f[521] && !f[304] && f[378];
	assign leaf[1692] = f[439] && f[521] && f[304] && !f[382];
	assign leaf[1693] = f[439] && f[521] && f[304] && f[382];
	
	// Tree 109, Classifier 9, Iteration: 10
	assign leaf[1694] = !f[568] && !f[720] && !f[177] && !f[294];
	assign leaf[1695] = !f[568] && !f[720] && !f[177] && f[294];
	assign leaf[1696] = !f[568] && !f[720] && f[177] && !f[287];
	assign leaf[1697] = !f[568] && !f[720] && f[177] && f[287];
	assign leaf[1698] = !f[568] && f[720] && !f[717] && !f[202];
	assign leaf[1699] = !f[568] && f[720] && !f[717] && f[202];
	assign leaf[1700] = !f[568] && f[720] && f[717] && !f[429];
	assign leaf[1701] = !f[568] && f[720] && f[717] && f[429];
	assign leaf[1702] = f[568] && !f[341] && !f[689] && !f[676];
	assign leaf[1703] = f[568] && !f[341] && !f[689] && f[676];
	assign leaf[1704] = f[568] && !f[341] && f[689] && !f[625];
	assign leaf[1705] = f[568] && !f[341] && f[689] && f[625];
	assign leaf[1706] = f[568] && f[341] && !f[543] && !f[573];
	assign leaf[1707] = f[568] && f[341] && !f[543] && f[573];
	assign leaf[1708] = f[568] && f[341] && f[543] && !f[576];
	assign leaf[1709] = f[568] && f[341] && f[543] && f[576];
	
	// Tree 110, Classifier 0, Iteration: 11
	assign leaf[1710] = !f[379] && !f[491] && !f[323] && !f[436];
	assign leaf[1711] = !f[379] && !f[491] && !f[323] && f[436];
	assign leaf[1712] = !f[379] && !f[491] && f[323] && !f[239];
	assign leaf[1713] = !f[379] && !f[491] && f[323] && f[239];
	assign leaf[1714] = !f[379] && f[491] && !f[348] && !f[387];
	assign leaf[1715] = !f[379] && f[491] && !f[348] && f[387];
	assign leaf[1716] = !f[379] && f[491] && f[348] && !f[625];
	assign leaf[1717] = !f[379] && f[491] && f[348] && f[625];
	assign leaf[1718] = f[379] && !f[329] && !f[331] && !f[513];
	assign leaf[1719] = f[379] && !f[329] && !f[331] && f[513];
	assign leaf[1720] = f[379] && !f[329] && f[331] && !f[346];
	assign leaf[1721] = f[379] && !f[329] && f[331] && f[346];
	assign leaf[1722] = f[379] && f[329] && !f[215] && !f[443];
	assign leaf[1723] = f[379] && f[329] && !f[215] && f[443];
	assign leaf[1724] = f[379] && f[329] && f[215] && !f[382];
	assign leaf[1725] = f[379] && f[329] && f[215] && f[382];
	
	// Tree 111, Classifier 1, Iteration: 11
	assign leaf[1726] = !f[466] && !f[374] && !f[511] && !f[683];
	assign leaf[1727] = !f[466] && !f[374] && !f[511] && f[683];
	assign leaf[1728] = !f[466] && !f[374] && f[511] && !f[649];
	assign leaf[1729] = !f[466] && !f[374] && f[511] && f[649];
	assign leaf[1730] = !f[466] && f[374] && !f[294];
	assign leaf[1731] = !f[466] && f[374] && f[294] && !f[404];
	assign leaf[1732] = !f[466] && f[374] && f[294] && f[404];
	assign leaf[1733] = f[466] && !f[145] && !f[556] && !f[467];
	assign leaf[1734] = f[466] && !f[145] && !f[556] && f[467];
	assign leaf[1735] = f[466] && !f[145] && f[556];
	assign leaf[1736] = f[466] && f[145];
	
	// Tree 112, Classifier 2, Iteration: 11
	assign leaf[1737] = !f[580] && !f[525] && !f[635] && !f[471];
	assign leaf[1738] = !f[580] && !f[525] && !f[635] && f[471];
	assign leaf[1739] = !f[580] && !f[525] && f[635] && !f[551];
	assign leaf[1740] = !f[580] && !f[525] && f[635] && f[551];
	assign leaf[1741] = !f[580] && f[525] && !f[605] && !f[387];
	assign leaf[1742] = !f[580] && f[525] && !f[605] && f[387];
	assign leaf[1743] = !f[580] && f[525] && f[605] && !f[434];
	assign leaf[1744] = !f[580] && f[525] && f[605] && f[434];
	assign leaf[1745] = f[580] && !f[468] && !f[414] && !f[662];
	assign leaf[1746] = f[580] && !f[468] && !f[414] && f[662];
	assign leaf[1747] = f[580] && !f[468] && f[414];
	assign leaf[1748] = f[580] && f[468] && !f[520] && !f[131];
	assign leaf[1749] = f[580] && f[468] && !f[520] && f[131];
	assign leaf[1750] = f[580] && f[468] && f[520] && !f[371];
	assign leaf[1751] = f[580] && f[468] && f[520] && f[371];
	
	// Tree 113, Classifier 3, Iteration: 11
	assign leaf[1752] = !f[428] && !f[523] && !f[565] && !f[181];
	assign leaf[1753] = !f[428] && !f[523] && !f[565] && f[181];
	assign leaf[1754] = !f[428] && !f[523] && f[565] && !f[353];
	assign leaf[1755] = !f[428] && !f[523] && f[565] && f[353];
	assign leaf[1756] = !f[428] && f[523] && !f[240] && !f[243];
	assign leaf[1757] = !f[428] && f[523] && !f[240] && f[243];
	assign leaf[1758] = !f[428] && f[523] && f[240] && !f[516];
	assign leaf[1759] = !f[428] && f[523] && f[240] && f[516];
	assign leaf[1760] = f[428] && !f[680] && !f[343] && !f[202];
	assign leaf[1761] = f[428] && !f[680] && !f[343] && f[202];
	assign leaf[1762] = f[428] && !f[680] && f[343] && !f[318];
	assign leaf[1763] = f[428] && !f[680] && f[343] && f[318];
	assign leaf[1764] = f[428] && f[680] && !f[318] && !f[539];
	assign leaf[1765] = f[428] && f[680] && !f[318] && f[539];
	assign leaf[1766] = f[428] && f[680] && f[318] && !f[204];
	assign leaf[1767] = f[428] && f[680] && f[318] && f[204];
	
	// Tree 114, Classifier 4, Iteration: 11
	assign leaf[1768] = !f[437] && !f[577] && !f[322] && !f[239];
	assign leaf[1769] = !f[437] && !f[577] && !f[322] && f[239];
	assign leaf[1770] = !f[437] && !f[577] && f[322] && !f[408];
	assign leaf[1771] = !f[437] && !f[577] && f[322] && f[408];
	assign leaf[1772] = !f[437] && f[577] && !f[690] && !f[438];
	assign leaf[1773] = !f[437] && f[577] && !f[690] && f[438];
	assign leaf[1774] = !f[437] && f[577] && f[690] && !f[269];
	assign leaf[1775] = !f[437] && f[577] && f[690] && f[269];
	assign leaf[1776] = f[437] && !f[461] && !f[434] && !f[484];
	assign leaf[1777] = f[437] && !f[461] && !f[434] && f[484];
	assign leaf[1778] = f[437] && !f[461] && f[434] && !f[598];
	assign leaf[1779] = f[437] && !f[461] && f[434] && f[598];
	assign leaf[1780] = f[437] && f[461] && !f[542] && !f[234];
	assign leaf[1781] = f[437] && f[461] && !f[542] && f[234];
	assign leaf[1782] = f[437] && f[461] && f[542] && !f[183];
	assign leaf[1783] = f[437] && f[461] && f[542] && f[183];
	
	// Tree 115, Classifier 5, Iteration: 11
	assign leaf[1784] = !f[190] && !f[248] && !f[491] && !f[268];
	assign leaf[1785] = !f[190] && !f[248] && !f[491] && f[268];
	assign leaf[1786] = !f[190] && !f[248] && f[491] && !f[304];
	assign leaf[1787] = !f[190] && !f[248] && f[491] && f[304];
	assign leaf[1788] = !f[190] && f[248] && !f[355] && !f[359];
	assign leaf[1789] = !f[190] && f[248] && !f[355] && f[359];
	assign leaf[1790] = !f[190] && f[248] && f[355] && !f[350];
	assign leaf[1791] = !f[190] && f[248] && f[355] && f[350];
	assign leaf[1792] = f[190] && !f[301] && !f[303] && !f[299];
	assign leaf[1793] = f[190] && !f[301] && !f[303] && f[299];
	assign leaf[1794] = f[190] && !f[301] && f[303] && !f[434];
	assign leaf[1795] = f[190] && !f[301] && f[303] && f[434];
	assign leaf[1796] = f[190] && f[301] && !f[269];
	assign leaf[1797] = f[190] && f[301] && f[269] && !f[329];
	assign leaf[1798] = f[190] && f[301] && f[269] && f[329];
	
	// Tree 116, Classifier 6, Iteration: 11
	assign leaf[1799] = !f[573] && !f[600] && !f[387] && !f[68];
	assign leaf[1800] = !f[573] && !f[600] && !f[387] && f[68];
	assign leaf[1801] = !f[573] && !f[600] && f[387] && !f[520];
	assign leaf[1802] = !f[573] && !f[600] && f[387] && f[520];
	assign leaf[1803] = !f[573] && f[600] && !f[458] && !f[427];
	assign leaf[1804] = !f[573] && f[600] && !f[458] && f[427];
	assign leaf[1805] = !f[573] && f[600] && f[458] && !f[297];
	assign leaf[1806] = !f[573] && f[600] && f[458] && f[297];
	assign leaf[1807] = f[573] && !f[656] && !f[625] && !f[240];
	assign leaf[1808] = f[573] && !f[656] && !f[625] && f[240];
	assign leaf[1809] = f[573] && !f[656] && f[625] && !f[107];
	assign leaf[1810] = f[573] && !f[656] && f[625] && f[107];
	assign leaf[1811] = f[573] && f[656] && !f[132] && !f[134];
	assign leaf[1812] = f[573] && f[656] && !f[132] && f[134];
	assign leaf[1813] = f[573] && f[656] && f[132] && !f[381];
	assign leaf[1814] = f[573] && f[656] && f[132] && f[381];
	
	// Tree 117, Classifier 7, Iteration: 11
	assign leaf[1815] = !f[376] && !f[297] && !f[707] && !f[232];
	assign leaf[1816] = !f[376] && !f[297] && !f[707] && f[232];
	assign leaf[1817] = !f[376] && !f[297] && f[707] && !f[243];
	assign leaf[1818] = !f[376] && !f[297] && f[707] && f[243];
	assign leaf[1819] = !f[376] && f[297] && !f[266] && !f[607];
	assign leaf[1820] = !f[376] && f[297] && !f[266] && f[607];
	assign leaf[1821] = !f[376] && f[297] && f[266] && !f[581];
	assign leaf[1822] = !f[376] && f[297] && f[266] && f[581];
	assign leaf[1823] = f[376] && !f[312] && !f[184] && !f[355];
	assign leaf[1824] = f[376] && !f[312] && !f[184] && f[355];
	assign leaf[1825] = f[376] && !f[312] && f[184] && !f[347];
	assign leaf[1826] = f[376] && !f[312] && f[184] && f[347];
	assign leaf[1827] = f[376] && f[312] && !f[581] && !f[346];
	assign leaf[1828] = f[376] && f[312] && !f[581] && f[346];
	assign leaf[1829] = f[376] && f[312] && f[581] && !f[413];
	assign leaf[1830] = f[376] && f[312] && f[581] && f[413];
	
	// Tree 118, Classifier 8, Iteration: 11
	assign leaf[1831] = !f[438] && !f[434] && !f[378] && !f[410];
	assign leaf[1832] = !f[438] && !f[434] && !f[378] && f[410];
	assign leaf[1833] = !f[438] && !f[434] && f[378] && !f[153];
	assign leaf[1834] = !f[438] && !f[434] && f[378] && f[153];
	assign leaf[1835] = !f[438] && f[434] && !f[687] && !f[292];
	assign leaf[1836] = !f[438] && f[434] && !f[687] && f[292];
	assign leaf[1837] = !f[438] && f[434] && f[687] && !f[544];
	assign leaf[1838] = !f[438] && f[434] && f[687] && f[544];
	assign leaf[1839] = f[438] && !f[520] && !f[330] && !f[153];
	assign leaf[1840] = f[438] && !f[520] && !f[330] && f[153];
	assign leaf[1841] = f[438] && !f[520] && f[330] && !f[300];
	assign leaf[1842] = f[438] && !f[520] && f[330] && f[300];
	assign leaf[1843] = f[438] && f[520] && !f[302] && !f[331];
	assign leaf[1844] = f[438] && f[520] && !f[302] && f[331];
	assign leaf[1845] = f[438] && f[520] && f[302] && !f[427];
	assign leaf[1846] = f[438] && f[520] && f[302] && f[427];
	
	// Tree 119, Classifier 9, Iteration: 11
	assign leaf[1847] = !f[158] && !f[126] && !f[218] && !f[400];
	assign leaf[1848] = !f[158] && !f[126] && !f[218] && f[400];
	assign leaf[1849] = !f[158] && !f[126] && f[218] && !f[214];
	assign leaf[1850] = !f[158] && !f[126] && f[218] && f[214];
	assign leaf[1851] = !f[158] && f[126] && !f[626];
	assign leaf[1852] = !f[158] && f[126] && f[626] && !f[261];
	assign leaf[1853] = !f[158] && f[126] && f[626] && f[261];
	assign leaf[1854] = f[158] && !f[329] && !f[518] && !f[356];
	assign leaf[1855] = f[158] && !f[329] && !f[518] && f[356];
	assign leaf[1856] = f[158] && !f[329] && f[518] && !f[241];
	assign leaf[1857] = f[158] && !f[329] && f[518] && f[241];
	assign leaf[1858] = f[158] && f[329] && !f[372] && !f[371];
	assign leaf[1859] = f[158] && f[329] && !f[372] && f[371];
	assign leaf[1860] = f[158] && f[329] && f[372] && !f[411];
	assign leaf[1861] = f[158] && f[329] && f[372] && f[411];
	
	// Tree 120, Classifier 0, Iteration: 12
	assign leaf[1862] = !f[387] && !f[429] && !f[427] && !f[430];
	assign leaf[1863] = !f[387] && !f[429] && !f[427] && f[430];
	assign leaf[1864] = !f[387] && !f[429] && f[427] && !f[625];
	assign leaf[1865] = !f[387] && !f[429] && f[427] && f[625];
	assign leaf[1866] = !f[387] && f[429] && !f[627] && !f[624];
	assign leaf[1867] = !f[387] && f[429] && !f[627] && f[624];
	assign leaf[1868] = !f[387] && f[429] && f[627] && !f[513];
	assign leaf[1869] = !f[387] && f[429] && f[627] && f[513];
	assign leaf[1870] = f[387] && !f[426] && !f[302] && !f[304];
	assign leaf[1871] = f[387] && !f[426] && !f[302] && f[304];
	assign leaf[1872] = f[387] && !f[426] && f[302] && !f[539];
	assign leaf[1873] = f[387] && !f[426] && f[302] && f[539];
	assign leaf[1874] = f[387] && f[426] && !f[437] && !f[433];
	assign leaf[1875] = f[387] && f[426] && !f[437] && f[433];
	assign leaf[1876] = f[387] && f[426] && f[437] && !f[301];
	assign leaf[1877] = f[387] && f[426] && f[437] && f[301];
	
	// Tree 121, Classifier 1, Iteration: 12
	assign leaf[1878] = !f[438] && !f[235] && !f[493] && !f[150];
	assign leaf[1879] = !f[438] && !f[235] && !f[493] && f[150];
	assign leaf[1880] = !f[438] && !f[235] && f[493] && !f[181];
	assign leaf[1881] = !f[438] && !f[235] && f[493] && f[181];
	assign leaf[1882] = !f[438] && f[235] && !f[151] && !f[98];
	assign leaf[1883] = !f[438] && f[235] && !f[151] && f[98];
	assign leaf[1884] = !f[438] && f[235] && f[151] && !f[265];
	assign leaf[1885] = !f[438] && f[235] && f[151] && f[265];
	assign leaf[1886] = f[438] && !f[439] && !f[609] && !f[123];
	assign leaf[1887] = f[438] && !f[439] && !f[609] && f[123];
	assign leaf[1888] = f[438] && !f[439] && f[609];
	assign leaf[1889] = f[438] && f[439] && !f[163];
	assign leaf[1890] = f[438] && f[439] && f[163];
	
	// Tree 122, Classifier 2, Iteration: 12
	assign leaf[1891] = !f[128] && !f[149] && !f[516] && !f[473];
	assign leaf[1892] = !f[128] && !f[149] && !f[516] && f[473];
	assign leaf[1893] = !f[128] && !f[149] && f[516] && !f[526];
	assign leaf[1894] = !f[128] && !f[149] && f[516] && f[526];
	assign leaf[1895] = !f[128] && f[149] && !f[317] && !f[259];
	assign leaf[1896] = !f[128] && f[149] && !f[317] && f[259];
	assign leaf[1897] = !f[128] && f[149] && f[317] && !f[155];
	assign leaf[1898] = !f[128] && f[149] && f[317] && f[155];
	assign leaf[1899] = f[128] && !f[630] && !f[294] && !f[292];
	assign leaf[1900] = f[128] && !f[630] && !f[294] && f[292];
	assign leaf[1901] = f[128] && !f[630] && f[294] && !f[607];
	assign leaf[1902] = f[128] && !f[630] && f[294] && f[607];
	assign leaf[1903] = f[128] && f[630] && !f[487] && !f[352];
	assign leaf[1904] = f[128] && f[630] && !f[487] && f[352];
	assign leaf[1905] = f[128] && f[630] && f[487] && !f[464];
	assign leaf[1906] = f[128] && f[630] && f[487] && f[464];
	
	// Tree 123, Classifier 3, Iteration: 12
	assign leaf[1907] = !f[371] && !f[291] && !f[182] && !f[578];
	assign leaf[1908] = !f[371] && !f[291] && !f[182] && f[578];
	assign leaf[1909] = !f[371] && !f[291] && f[182] && !f[317];
	assign leaf[1910] = !f[371] && !f[291] && f[182] && f[317];
	assign leaf[1911] = !f[371] && f[291] && !f[266] && !f[651];
	assign leaf[1912] = !f[371] && f[291] && !f[266] && f[651];
	assign leaf[1913] = !f[371] && f[291] && f[266] && !f[123];
	assign leaf[1914] = !f[371] && f[291] && f[266] && f[123];
	assign leaf[1915] = f[371] && !f[320] && !f[259] && !f[149];
	assign leaf[1916] = f[371] && !f[320] && !f[259] && f[149];
	assign leaf[1917] = f[371] && !f[320] && f[259] && !f[375];
	assign leaf[1918] = f[371] && !f[320] && f[259] && f[375];
	assign leaf[1919] = f[371] && f[320] && !f[151] && !f[256];
	assign leaf[1920] = f[371] && f[320] && !f[151] && f[256];
	assign leaf[1921] = f[371] && f[320] && f[151] && !f[260];
	assign leaf[1922] = f[371] && f[320] && f[151] && f[260];
	
	// Tree 124, Classifier 4, Iteration: 12
	assign leaf[1923] = !f[346] && !f[208] && !f[465] && !f[637];
	assign leaf[1924] = !f[346] && !f[208] && !f[465] && f[637];
	assign leaf[1925] = !f[346] && !f[208] && f[465] && !f[291];
	assign leaf[1926] = !f[346] && !f[208] && f[465] && f[291];
	assign leaf[1927] = !f[346] && f[208] && !f[211] && !f[218];
	assign leaf[1928] = !f[346] && f[208] && !f[211] && f[218];
	assign leaf[1929] = !f[346] && f[208] && f[211] && !f[248];
	assign leaf[1930] = !f[346] && f[208] && f[211] && f[248];
	assign leaf[1931] = f[346] && !f[427] && !f[551] && !f[238];
	assign leaf[1932] = f[346] && !f[427] && !f[551] && f[238];
	assign leaf[1933] = f[346] && !f[427] && f[551] && !f[603];
	assign leaf[1934] = f[346] && !f[427] && f[551] && f[603];
	assign leaf[1935] = f[346] && f[427] && !f[568] && !f[710];
	assign leaf[1936] = f[346] && f[427] && !f[568] && f[710];
	assign leaf[1937] = f[346] && f[427] && f[568] && !f[157];
	assign leaf[1938] = f[346] && f[427] && f[568] && f[157];
	
	// Tree 125, Classifier 5, Iteration: 12
	assign leaf[1939] = !f[485] && !f[160] && !f[218] && !f[435];
	assign leaf[1940] = !f[485] && !f[160] && !f[218] && f[435];
	assign leaf[1941] = !f[485] && !f[160] && f[218] && !f[331];
	assign leaf[1942] = !f[485] && !f[160] && f[218] && f[331];
	assign leaf[1943] = !f[485] && f[160] && !f[271] && !f[246];
	assign leaf[1944] = !f[485] && f[160] && !f[271] && f[246];
	assign leaf[1945] = !f[485] && f[160] && f[271] && !f[687];
	assign leaf[1946] = !f[485] && f[160] && f[271] && f[687];
	assign leaf[1947] = f[485] && !f[458] && !f[428] && !f[349];
	assign leaf[1948] = f[485] && !f[458] && !f[428] && f[349];
	assign leaf[1949] = f[485] && !f[458] && f[428] && !f[512];
	assign leaf[1950] = f[485] && !f[458] && f[428] && f[512];
	assign leaf[1951] = f[485] && f[458] && !f[513] && !f[355];
	assign leaf[1952] = f[485] && f[458] && !f[513] && f[355];
	assign leaf[1953] = f[485] && f[458] && f[513] && !f[177];
	assign leaf[1954] = f[485] && f[458] && f[513] && f[177];
	
	// Tree 126, Classifier 6, Iteration: 12
	assign leaf[1955] = !f[269] && !f[654] && !f[576] && !f[548];
	assign leaf[1956] = !f[269] && !f[654] && !f[576] && f[548];
	assign leaf[1957] = !f[269] && !f[654] && f[576] && !f[660];
	assign leaf[1958] = !f[269] && !f[654] && f[576] && f[660];
	assign leaf[1959] = !f[269] && f[654] && !f[134] && !f[131];
	assign leaf[1960] = !f[269] && f[654] && !f[134] && f[131];
	assign leaf[1961] = !f[269] && f[654] && f[134] && !f[353];
	assign leaf[1962] = !f[269] && f[654] && f[134] && f[353];
	assign leaf[1963] = f[269] && !f[163] && !f[357] && !f[132];
	assign leaf[1964] = f[269] && !f[163] && !f[357] && f[132];
	assign leaf[1965] = f[269] && !f[163] && f[357] && !f[239];
	assign leaf[1966] = f[269] && !f[163] && f[357] && f[239];
	assign leaf[1967] = f[269] && f[163] && !f[349];
	assign leaf[1968] = f[269] && f[163] && f[349] && !f[622];
	assign leaf[1969] = f[269] && f[163] && f[349] && f[622];
	
	// Tree 127, Classifier 7, Iteration: 12
	assign leaf[1970] = !f[158] && !f[153] && !f[432] && !f[377];
	assign leaf[1971] = !f[158] && !f[153] && !f[432] && f[377];
	assign leaf[1972] = !f[158] && !f[153] && f[432] && !f[372];
	assign leaf[1973] = !f[158] && !f[153] && f[432] && f[372];
	assign leaf[1974] = !f[158] && f[153] && !f[604] && !f[634];
	assign leaf[1975] = !f[158] && f[153] && !f[604] && f[634];
	assign leaf[1976] = !f[158] && f[153] && f[604] && !f[687];
	assign leaf[1977] = !f[158] && f[153] && f[604] && f[687];
	assign leaf[1978] = f[158] && !f[686] && !f[149] && !f[687];
	assign leaf[1979] = f[158] && !f[686] && !f[149] && f[687];
	assign leaf[1980] = f[158] && !f[686] && f[149] && !f[605];
	assign leaf[1981] = f[158] && !f[686] && f[149] && f[605];
	assign leaf[1982] = f[158] && f[686] && !f[573];
	assign leaf[1983] = f[158] && f[686] && f[573] && !f[374];
	assign leaf[1984] = f[158] && f[686] && f[573] && f[374];
	
	// Tree 128, Classifier 8, Iteration: 12
	assign leaf[1985] = !f[274] && !f[660] && !f[597] && !f[567];
	assign leaf[1986] = !f[274] && !f[660] && !f[597] && f[567];
	assign leaf[1987] = !f[274] && !f[660] && f[597] && !f[572];
	assign leaf[1988] = !f[274] && !f[660] && f[597] && f[572];
	assign leaf[1989] = !f[274] && f[660] && !f[544] && !f[542];
	assign leaf[1990] = !f[274] && f[660] && !f[544] && f[542];
	assign leaf[1991] = !f[274] && f[660] && f[544] && !f[513];
	assign leaf[1992] = !f[274] && f[660] && f[544] && f[513];
	assign leaf[1993] = f[274] && !f[426] && !f[271] && !f[380];
	assign leaf[1994] = f[274] && !f[426] && !f[271] && f[380];
	assign leaf[1995] = f[274] && !f[426] && f[271] && !f[486];
	assign leaf[1996] = f[274] && !f[426] && f[271] && f[486];
	assign leaf[1997] = f[274] && f[426] && !f[520] && !f[409];
	assign leaf[1998] = f[274] && f[426] && !f[520] && f[409];
	assign leaf[1999] = f[274] && f[426] && f[520] && !f[634];
	assign leaf[2000] = f[274] && f[426] && f[520] && f[634];
	
	// Tree 129, Classifier 9, Iteration: 12
	assign leaf[2001] = !f[719] && !f[578] && !f[318] && !f[316];
	assign leaf[2002] = !f[719] && !f[578] && !f[318] && f[316];
	assign leaf[2003] = !f[719] && !f[578] && f[318] && !f[468];
	assign leaf[2004] = !f[719] && !f[578] && f[318] && f[468];
	assign leaf[2005] = !f[719] && f[578] && !f[399] && !f[718];
	assign leaf[2006] = !f[719] && f[578] && !f[399] && f[718];
	assign leaf[2007] = !f[719] && f[578] && f[399] && !f[346];
	assign leaf[2008] = !f[719] && f[578] && f[399] && f[346];
	assign leaf[2009] = f[719] && !f[717] && !f[201] && !f[319];
	assign leaf[2010] = f[719] && !f[717] && !f[201] && f[319];
	assign leaf[2011] = f[719] && !f[717] && f[201] && !f[459];
	assign leaf[2012] = f[719] && !f[717] && f[201] && f[459];
	assign leaf[2013] = f[719] && f[717] && !f[431] && !f[458];
	assign leaf[2014] = f[719] && f[717] && !f[431] && f[458];
	assign leaf[2015] = f[719] && f[717] && f[431] && !f[633];
	assign leaf[2016] = f[719] && f[717] && f[431] && f[633];
	
	// Tree 130, Classifier 0, Iteration: 13
	assign leaf[2017] = !f[434] && !f[242] && !f[387] && !f[240];
	assign leaf[2018] = !f[434] && !f[242] && !f[387] && f[240];
	assign leaf[2019] = !f[434] && !f[242] && f[387] && !f[350];
	assign leaf[2020] = !f[434] && !f[242] && f[387] && f[350];
	assign leaf[2021] = !f[434] && f[242] && !f[570] && !f[624];
	assign leaf[2022] = !f[434] && f[242] && !f[570] && f[624];
	assign leaf[2023] = !f[434] && f[242] && f[570] && !f[401];
	assign leaf[2024] = !f[434] && f[242] && f[570] && f[401];
	assign leaf[2025] = f[434] && !f[540] && !f[537];
	assign leaf[2026] = f[434] && !f[540] && f[537] && !f[323];
	assign leaf[2027] = f[434] && !f[540] && f[537] && f[323];
	assign leaf[2028] = f[434] && f[540] && !f[344] && !f[374];
	assign leaf[2029] = f[434] && f[540] && !f[344] && f[374];
	assign leaf[2030] = f[434] && f[540] && f[344] && !f[656];
	assign leaf[2031] = f[434] && f[540] && f[344] && f[656];
	
	// Tree 131, Classifier 1, Iteration: 13
	assign leaf[2032] = !f[429] && !f[354] && !f[272] && !f[462];
	assign leaf[2033] = !f[429] && !f[354] && !f[272] && f[462];
	assign leaf[2034] = !f[429] && !f[354] && f[272] && !f[518];
	assign leaf[2035] = !f[429] && !f[354] && f[272] && f[518];
	assign leaf[2036] = !f[429] && f[354] && !f[162] && !f[296];
	assign leaf[2037] = !f[429] && f[354] && !f[162] && f[296];
	assign leaf[2038] = !f[429] && f[354] && f[162] && !f[211];
	assign leaf[2039] = !f[429] && f[354] && f[162] && f[211];
	assign leaf[2040] = f[429] && !f[375];
	assign leaf[2041] = f[429] && f[375] && !f[687] && !f[679];
	assign leaf[2042] = f[429] && f[375] && !f[687] && f[679];
	assign leaf[2043] = f[429] && f[375] && f[687] && !f[345];
	assign leaf[2044] = f[429] && f[375] && f[687] && f[345];
	
	// Tree 132, Classifier 2, Iteration: 13
	assign leaf[2045] = !f[345] && !f[348] && !f[370] && !f[607];
	assign leaf[2046] = !f[345] && !f[348] && !f[370] && f[607];
	assign leaf[2047] = !f[345] && !f[348] && f[370] && !f[342];
	assign leaf[2048] = !f[345] && !f[348] && f[370] && f[342];
	assign leaf[2049] = !f[345] && f[348] && !f[581] && !f[526];
	assign leaf[2050] = !f[345] && f[348] && !f[581] && f[526];
	assign leaf[2051] = !f[345] && f[348] && f[581] && !f[440];
	assign leaf[2052] = !f[345] && f[348] && f[581] && f[440];
	assign leaf[2053] = f[345] && !f[401] && !f[515] && !f[186];
	assign leaf[2054] = f[345] && !f[401] && !f[515] && f[186];
	assign leaf[2055] = f[345] && !f[401] && f[515] && !f[293];
	assign leaf[2056] = f[345] && !f[401] && f[515] && f[293];
	assign leaf[2057] = f[345] && f[401] && !f[317] && !f[292];
	assign leaf[2058] = f[345] && f[401] && !f[317] && f[292];
	assign leaf[2059] = f[345] && f[401] && f[317] && !f[667];
	assign leaf[2060] = f[345] && f[401] && f[317] && f[667];
	
	// Tree 133, Classifier 3, Iteration: 13
	assign leaf[2061] = !f[456] && !f[518] && !f[515] && !f[342];
	assign leaf[2062] = !f[456] && !f[518] && !f[515] && f[342];
	assign leaf[2063] = !f[456] && !f[518] && f[515] && !f[460];
	assign leaf[2064] = !f[456] && !f[518] && f[515] && f[460];
	assign leaf[2065] = !f[456] && f[518] && !f[594] && !f[463];
	assign leaf[2066] = !f[456] && f[518] && !f[594] && f[463];
	assign leaf[2067] = !f[456] && f[518] && f[594] && !f[325];
	assign leaf[2068] = !f[456] && f[518] && f[594] && f[325];
	assign leaf[2069] = f[456] && !f[678] && !f[351] && !f[633];
	assign leaf[2070] = f[456] && !f[678] && !f[351] && f[633];
	assign leaf[2071] = f[456] && !f[678] && f[351] && !f[343];
	assign leaf[2072] = f[456] && !f[678] && f[351] && f[343];
	assign leaf[2073] = f[456] && f[678] && !f[292] && !f[322];
	assign leaf[2074] = f[456] && f[678] && !f[292] && f[322];
	assign leaf[2075] = f[456] && f[678] && f[292];
	
	// Tree 134, Classifier 4, Iteration: 13
	assign leaf[2076] = !f[595] && !f[374] && !f[426] && !f[373];
	assign leaf[2077] = !f[595] && !f[374] && !f[426] && f[373];
	assign leaf[2078] = !f[595] && !f[374] && f[426] && !f[294];
	assign leaf[2079] = !f[595] && !f[374] && f[426] && f[294];
	assign leaf[2080] = !f[595] && f[374] && !f[552] && !f[712];
	assign leaf[2081] = !f[595] && f[374] && !f[552] && f[712];
	assign leaf[2082] = !f[595] && f[374] && f[552] && !f[454];
	assign leaf[2083] = !f[595] && f[374] && f[552] && f[454];
	assign leaf[2084] = f[595] && !f[542] && !f[664];
	assign leaf[2085] = f[595] && !f[542] && f[664];
	assign leaf[2086] = f[595] && f[542] && !f[401] && !f[442];
	assign leaf[2087] = f[595] && f[542] && !f[401] && f[442];
	assign leaf[2088] = f[595] && f[542] && f[401] && !f[567];
	assign leaf[2089] = f[595] && f[542] && f[401] && f[567];
	
	// Tree 135, Classifier 5, Iteration: 13
	assign leaf[2090] = !f[346] && !f[459] && !f[568] && !f[189];
	assign leaf[2091] = !f[346] && !f[459] && !f[568] && f[189];
	assign leaf[2092] = !f[346] && !f[459] && f[568] && !f[293];
	assign leaf[2093] = !f[346] && !f[459] && f[568] && f[293];
	assign leaf[2094] = !f[346] && f[459] && !f[276] && !f[325];
	assign leaf[2095] = !f[346] && f[459] && !f[276] && f[325];
	assign leaf[2096] = !f[346] && f[459] && f[276] && !f[380];
	assign leaf[2097] = !f[346] && f[459] && f[276] && f[380];
	assign leaf[2098] = f[346] && !f[206] && !f[381] && !f[439];
	assign leaf[2099] = f[346] && !f[206] && !f[381] && f[439];
	assign leaf[2100] = f[346] && !f[206] && f[381] && !f[463];
	assign leaf[2101] = f[346] && !f[206] && f[381] && f[463];
	assign leaf[2102] = f[346] && f[206] && !f[269] && !f[266];
	assign leaf[2103] = f[346] && f[206] && !f[269] && f[266];
	assign leaf[2104] = f[346] && f[206] && f[269] && !f[238];
	assign leaf[2105] = f[346] && f[206] && f[269] && f[238];
	
	// Tree 136, Classifier 6, Iteration: 13
	assign leaf[2106] = !f[654] && !f[572] && !f[544] && !f[599];
	assign leaf[2107] = !f[654] && !f[572] && !f[544] && f[599];
	assign leaf[2108] = !f[654] && !f[572] && f[544] && !f[543];
	assign leaf[2109] = !f[654] && !f[572] && f[544] && f[543];
	assign leaf[2110] = !f[654] && f[572] && !f[429] && !f[431];
	assign leaf[2111] = !f[654] && f[572] && !f[429] && f[431];
	assign leaf[2112] = !f[654] && f[572] && f[429] && !f[593];
	assign leaf[2113] = !f[654] && f[572] && f[429] && f[593];
	assign leaf[2114] = f[654] && !f[132] && !f[131] && !f[164];
	assign leaf[2115] = f[654] && !f[132] && !f[131] && f[164];
	assign leaf[2116] = f[654] && !f[132] && f[131] && !f[430];
	assign leaf[2117] = f[654] && !f[132] && f[131] && f[430];
	assign leaf[2118] = f[654] && f[132] && !f[458] && !f[525];
	assign leaf[2119] = f[654] && f[132] && !f[458] && f[525];
	assign leaf[2120] = f[654] && f[132] && f[458] && !f[326];
	assign leaf[2121] = f[654] && f[132] && f[458] && f[326];
	
	// Tree 137, Classifier 7, Iteration: 13
	assign leaf[2122] = !f[569] && !f[267] && !f[433] && !f[487];
	assign leaf[2123] = !f[569] && !f[267] && !f[433] && f[487];
	assign leaf[2124] = !f[569] && !f[267] && f[433] && !f[346];
	assign leaf[2125] = !f[569] && !f[267] && f[433] && f[346];
	assign leaf[2126] = !f[569] && f[267] && !f[263] && !f[236];
	assign leaf[2127] = !f[569] && f[267] && !f[263] && f[236];
	assign leaf[2128] = !f[569] && f[267] && f[263] && !f[260];
	assign leaf[2129] = !f[569] && f[267] && f[263] && f[260];
	assign leaf[2130] = f[569] && !f[679] && !f[677] && !f[709];
	assign leaf[2131] = f[569] && !f[679] && !f[677] && f[709];
	assign leaf[2132] = f[569] && !f[679] && f[677] && !f[238];
	assign leaf[2133] = f[569] && !f[679] && f[677] && f[238];
	assign leaf[2134] = f[569] && f[679] && !f[271] && !f[326];
	assign leaf[2135] = f[569] && f[679] && !f[271] && f[326];
	assign leaf[2136] = f[569] && f[679] && f[271] && !f[602];
	assign leaf[2137] = f[569] && f[679] && f[271] && f[602];
	
	// Tree 138, Classifier 8, Iteration: 13
	assign leaf[2138] = !f[440] && !f[288] && !f[541] && !f[511];
	assign leaf[2139] = !f[440] && !f[288] && !f[541] && f[511];
	assign leaf[2140] = !f[440] && !f[288] && f[541] && !f[571];
	assign leaf[2141] = !f[440] && !f[288] && f[541] && f[571];
	assign leaf[2142] = !f[440] && f[288] && !f[374] && !f[348];
	assign leaf[2143] = !f[440] && f[288] && !f[374] && f[348];
	assign leaf[2144] = !f[440] && f[288] && f[374] && !f[517];
	assign leaf[2145] = !f[440] && f[288] && f[374] && f[517];
	assign leaf[2146] = f[440] && !f[582] && !f[304] && !f[494];
	assign leaf[2147] = f[440] && !f[582] && !f[304] && f[494];
	assign leaf[2148] = f[440] && !f[582] && f[304] && !f[371];
	assign leaf[2149] = f[440] && !f[582] && f[304] && f[371];
	assign leaf[2150] = f[440] && f[582] && !f[525] && !f[349];
	assign leaf[2151] = f[440] && f[582] && !f[525] && f[349];
	assign leaf[2152] = f[440] && f[582] && f[525] && !f[460];
	assign leaf[2153] = f[440] && f[582] && f[525] && f[460];
	
	// Tree 139, Classifier 9, Iteration: 13
	assign leaf[2154] = !f[159] && !f[632] && !f[212] && !f[572];
	assign leaf[2155] = !f[159] && !f[632] && !f[212] && f[572];
	assign leaf[2156] = !f[159] && !f[632] && f[212] && !f[291];
	assign leaf[2157] = !f[159] && !f[632] && f[212] && f[291];
	assign leaf[2158] = !f[159] && f[632] && !f[601] && !f[683];
	assign leaf[2159] = !f[159] && f[632] && !f[601] && f[683];
	assign leaf[2160] = !f[159] && f[632] && f[601] && !f[517];
	assign leaf[2161] = !f[159] && f[632] && f[601] && f[517];
	assign leaf[2162] = f[159] && !f[355] && !f[657] && !f[688];
	assign leaf[2163] = f[159] && !f[355] && !f[657] && f[688];
	assign leaf[2164] = f[159] && !f[355] && f[657];
	assign leaf[2165] = f[159] && f[355] && !f[290] && !f[682];
	assign leaf[2166] = f[159] && f[355] && !f[290] && f[682];
	assign leaf[2167] = f[159] && f[355] && f[290] && !f[493];
	assign leaf[2168] = f[159] && f[355] && f[290] && f[493];
	
	// Tree 140, Classifier 0, Iteration: 14
	assign leaf[2169] = !f[406] && !f[490] && !f[323] && !f[629];
	assign leaf[2170] = !f[406] && !f[490] && !f[323] && f[629];
	assign leaf[2171] = !f[406] && !f[490] && f[323] && !f[239];
	assign leaf[2172] = !f[406] && !f[490] && f[323] && f[239];
	assign leaf[2173] = !f[406] && f[490] && !f[294] && !f[415];
	assign leaf[2174] = !f[406] && f[490] && !f[294] && f[415];
	assign leaf[2175] = !f[406] && f[490] && f[294] && !f[570];
	assign leaf[2176] = !f[406] && f[490] && f[294] && f[570];
	assign leaf[2177] = f[406] && !f[329] && !f[332] && !f[328];
	assign leaf[2178] = f[406] && !f[329] && !f[332] && f[328];
	assign leaf[2179] = f[406] && !f[329] && f[332] && !f[656];
	assign leaf[2180] = f[406] && !f[329] && f[332] && f[656];
	assign leaf[2181] = f[406] && f[329] && !f[295] && !f[404];
	assign leaf[2182] = f[406] && f[329] && !f[295] && f[404];
	assign leaf[2183] = f[406] && f[329] && f[295] && !f[412];
	assign leaf[2184] = f[406] && f[329] && f[295] && f[412];
	
	// Tree 141, Classifier 1, Iteration: 14
	assign leaf[2185] = !f[355] && !f[684] && !f[467] && !f[510];
	assign leaf[2186] = !f[355] && !f[684] && !f[467] && f[510];
	assign leaf[2187] = !f[355] && !f[684] && f[467] && !f[98];
	assign leaf[2188] = !f[355] && !f[684] && f[467] && f[98];
	assign leaf[2189] = !f[355] && f[684] && !f[208] && !f[295];
	assign leaf[2190] = !f[355] && f[684] && !f[208] && f[295];
	assign leaf[2191] = !f[355] && f[684] && f[208] && !f[409];
	assign leaf[2192] = !f[355] && f[684] && f[208] && f[409];
	assign leaf[2193] = f[355] && !f[161] && !f[192] && !f[102];
	assign leaf[2194] = f[355] && !f[161] && !f[192] && f[102];
	assign leaf[2195] = f[355] && !f[161] && f[192];
	assign leaf[2196] = f[355] && f[161] && !f[211] && !f[651];
	assign leaf[2197] = f[355] && f[161] && !f[211] && f[651];
	assign leaf[2198] = f[355] && f[161] && f[211] && !f[659];
	assign leaf[2199] = f[355] && f[161] && f[211] && f[659];
	
	// Tree 142, Classifier 2, Iteration: 14
	assign leaf[2200] = !f[683] && !f[659] && !f[492] && !f[576];
	assign leaf[2201] = !f[683] && !f[659] && !f[492] && f[576];
	assign leaf[2202] = !f[683] && !f[659] && f[492] && !f[352];
	assign leaf[2203] = !f[683] && !f[659] && f[492] && f[352];
	assign leaf[2204] = !f[683] && f[659] && !f[544] && !f[514];
	assign leaf[2205] = !f[683] && f[659] && !f[544] && f[514];
	assign leaf[2206] = !f[683] && f[659] && f[544] && !f[494];
	assign leaf[2207] = !f[683] && f[659] && f[544] && f[494];
	assign leaf[2208] = f[683] && !f[403] && !f[691] && !f[598];
	assign leaf[2209] = f[683] && !f[403] && !f[691] && f[598];
	assign leaf[2210] = f[683] && !f[403] && f[691];
	assign leaf[2211] = f[683] && f[403] && !f[610];
	assign leaf[2212] = f[683] && f[403] && f[610] && !f[325];
	assign leaf[2213] = f[683] && f[403] && f[610] && f[325];
	
	// Tree 143, Classifier 3, Iteration: 14
	assign leaf[2214] = !f[351] && !f[546] && !f[294] && !f[682];
	assign leaf[2215] = !f[351] && !f[546] && !f[294] && f[682];
	assign leaf[2216] = !f[351] && !f[546] && f[294] && !f[298];
	assign leaf[2217] = !f[351] && !f[546] && f[294] && f[298];
	assign leaf[2218] = !f[351] && f[546] && !f[464] && !f[353];
	assign leaf[2219] = !f[351] && f[546] && !f[464] && f[353];
	assign leaf[2220] = !f[351] && f[546] && f[464] && !f[678];
	assign leaf[2221] = !f[351] && f[546] && f[464] && f[678];
	assign leaf[2222] = f[351] && !f[269] && !f[271] && !f[175];
	assign leaf[2223] = f[351] && !f[269] && !f[271] && f[175];
	assign leaf[2224] = f[351] && !f[269] && f[271] && !f[345];
	assign leaf[2225] = f[351] && !f[269] && f[271] && f[345];
	assign leaf[2226] = f[351] && f[269] && !f[183] && !f[127];
	assign leaf[2227] = f[351] && f[269] && !f[183] && f[127];
	assign leaf[2228] = f[351] && f[269] && f[183] && !f[514];
	assign leaf[2229] = f[351] && f[269] && f[183] && f[514];
	
	// Tree 144, Classifier 4, Iteration: 14
	assign leaf[2230] = !f[408] && !f[466] && !f[146] && !f[381];
	assign leaf[2231] = !f[408] && !f[466] && !f[146] && f[381];
	assign leaf[2232] = !f[408] && !f[466] && f[146];
	assign leaf[2233] = !f[408] && f[466] && !f[488] && !f[295];
	assign leaf[2234] = !f[408] && f[466] && !f[488] && f[295];
	assign leaf[2235] = !f[408] && f[466] && f[488] && !f[572];
	assign leaf[2236] = !f[408] && f[466] && f[488] && f[572];
	assign leaf[2237] = f[408] && !f[209] && !f[544] && !f[627];
	assign leaf[2238] = f[408] && !f[209] && !f[544] && f[627];
	assign leaf[2239] = f[408] && !f[209] && f[544] && !f[551];
	assign leaf[2240] = f[408] && !f[209] && f[544] && f[551];
	assign leaf[2241] = f[408] && f[209] && !f[212] && !f[205];
	assign leaf[2242] = f[408] && f[209] && !f[212] && f[205];
	assign leaf[2243] = f[408] && f[209] && f[212] && !f[320];
	assign leaf[2244] = f[408] && f[209] && f[212] && f[320];
	
	// Tree 145, Classifier 5, Iteration: 14
	assign leaf[2245] = !f[488] && !f[457] && !f[159] && !f[217];
	assign leaf[2246] = !f[488] && !f[457] && !f[159] && f[217];
	assign leaf[2247] = !f[488] && !f[457] && f[159] && !f[271];
	assign leaf[2248] = !f[488] && !f[457] && f[159] && f[271];
	assign leaf[2249] = !f[488] && f[457] && !f[513] && !f[483];
	assign leaf[2250] = !f[488] && f[457] && !f[513] && f[483];
	assign leaf[2251] = !f[488] && f[457] && f[513] && !f[430];
	assign leaf[2252] = !f[488] && f[457] && f[513] && f[430];
	assign leaf[2253] = f[488] && !f[380] && !f[686] && !f[276];
	assign leaf[2254] = f[488] && !f[380] && !f[686] && f[276];
	assign leaf[2255] = f[488] && !f[380] && f[686] && !f[378];
	assign leaf[2256] = f[488] && !f[380] && f[686] && f[378];
	assign leaf[2257] = f[488] && f[380] && !f[434] && !f[540];
	assign leaf[2258] = f[488] && f[380] && !f[434] && f[540];
	assign leaf[2259] = f[488] && f[380] && f[434] && !f[551];
	assign leaf[2260] = f[488] && f[380] && f[434] && f[551];
	
	// Tree 146, Classifier 6, Iteration: 14
	assign leaf[2261] = !f[242] && !f[296] && !f[216] && !f[350];
	assign leaf[2262] = !f[242] && !f[296] && !f[216] && f[350];
	assign leaf[2263] = !f[242] && !f[296] && f[216] && !f[632];
	assign leaf[2264] = !f[242] && !f[296] && f[216] && f[632];
	assign leaf[2265] = !f[242] && f[296] && !f[357] && !f[131];
	assign leaf[2266] = !f[242] && f[296] && !f[357] && f[131];
	assign leaf[2267] = !f[242] && f[296] && f[357] && !f[485];
	assign leaf[2268] = !f[242] && f[296] && f[357] && f[485];
	assign leaf[2269] = f[242] && !f[164] && !f[326] && !f[131];
	assign leaf[2270] = f[242] && !f[164] && !f[326] && f[131];
	assign leaf[2271] = f[242] && !f[164] && f[326] && !f[387];
	assign leaf[2272] = f[242] && !f[164] && f[326] && f[387];
	assign leaf[2273] = f[242] && f[164] && !f[623];
	assign leaf[2274] = f[242] && f[164] && f[623] && !f[622];
	assign leaf[2275] = f[242] && f[164] && f[623] && f[622];
	
	// Tree 147, Classifier 7, Iteration: 14
	assign leaf[2276] = !f[580] && !f[259] && !f[206] && !f[459];
	assign leaf[2277] = !f[580] && !f[259] && !f[206] && f[459];
	assign leaf[2278] = !f[580] && !f[259] && f[206] && !f[578];
	assign leaf[2279] = !f[580] && !f[259] && f[206] && f[578];
	assign leaf[2280] = !f[580] && f[259] && !f[263] && !f[427];
	assign leaf[2281] = !f[580] && f[259] && !f[263] && f[427];
	assign leaf[2282] = !f[580] && f[259] && f[263] && !f[554];
	assign leaf[2283] = !f[580] && f[259] && f[263] && f[554];
	assign leaf[2284] = f[580] && !f[746] && !f[283] && !f[749];
	assign leaf[2285] = f[580] && !f[746] && !f[283] && f[749];
	assign leaf[2286] = f[580] && !f[746] && f[283] && !f[206];
	assign leaf[2287] = f[580] && !f[746] && f[283] && f[206];
	assign leaf[2288] = f[580] && f[746] && !f[436];
	assign leaf[2289] = f[580] && f[746] && f[436];
	
	// Tree 148, Classifier 8, Iteration: 14
	assign leaf[2290] = !f[466] && !f[185] && !f[157] && !f[627];
	assign leaf[2291] = !f[466] && !f[185] && !f[157] && f[627];
	assign leaf[2292] = !f[466] && !f[185] && f[157] && !f[580];
	assign leaf[2293] = !f[466] && !f[185] && f[157] && f[580];
	assign leaf[2294] = !f[466] && f[185] && !f[268] && !f[322];
	assign leaf[2295] = !f[466] && f[185] && !f[268] && f[322];
	assign leaf[2296] = !f[466] && f[185] && f[268] && !f[659];
	assign leaf[2297] = !f[466] && f[185] && f[268] && f[659];
	assign leaf[2298] = f[466] && !f[520] && !f[350] && !f[233];
	assign leaf[2299] = f[466] && !f[520] && !f[350] && f[233];
	assign leaf[2300] = f[466] && !f[520] && f[350] && !f[440];
	assign leaf[2301] = f[466] && !f[520] && f[350] && f[440];
	assign leaf[2302] = f[466] && f[520] && !f[180] && !f[620];
	assign leaf[2303] = f[466] && f[520] && !f[180] && f[620];
	assign leaf[2304] = f[466] && f[520] && f[180] && !f[275];
	assign leaf[2305] = f[466] && f[520] && f[180] && f[275];
	
	// Tree 149, Classifier 9, Iteration: 14
	assign leaf[2306] = !f[469] && !f[436] && !f[438] && !f[468];
	assign leaf[2307] = !f[469] && !f[436] && !f[438] && f[468];
	assign leaf[2308] = !f[469] && !f[436] && f[438] && !f[320];
	assign leaf[2309] = !f[469] && !f[436] && f[438] && f[320];
	assign leaf[2310] = !f[469] && f[436] && !f[567] && !f[233];
	assign leaf[2311] = !f[469] && f[436] && !f[567] && f[233];
	assign leaf[2312] = !f[469] && f[436] && f[567] && !f[398];
	assign leaf[2313] = !f[469] && f[436] && f[567] && f[398];
	assign leaf[2314] = f[469] && !f[369] && !f[694] && !f[385];
	assign leaf[2315] = f[469] && !f[369] && !f[694] && f[385];
	assign leaf[2316] = f[469] && !f[369] && f[694];
	assign leaf[2317] = f[469] && f[369] && !f[385] && !f[667];
	assign leaf[2318] = f[469] && f[369] && !f[385] && f[667];
	assign leaf[2319] = f[469] && f[369] && f[385] && !f[229];
	assign leaf[2320] = f[469] && f[369] && f[385] && f[229];
	
	// Tree 150, Classifier 0, Iteration: 15
	assign leaf[2321] = !f[379] && !f[491] && !f[322] && !f[435];
	assign leaf[2322] = !f[379] && !f[491] && !f[322] && f[435];
	assign leaf[2323] = !f[379] && !f[491] && f[322] && !f[273];
	assign leaf[2324] = !f[379] && !f[491] && f[322] && f[273];
	assign leaf[2325] = !f[379] && f[491] && !f[348] && !f[415];
	assign leaf[2326] = !f[379] && f[491] && !f[348] && f[415];
	assign leaf[2327] = !f[379] && f[491] && f[348] && !f[598];
	assign leaf[2328] = !f[379] && f[491] && f[348] && f[598];
	assign leaf[2329] = f[379] && !f[329] && !f[331] && !f[486];
	assign leaf[2330] = f[379] && !f[329] && !f[331] && f[486];
	assign leaf[2331] = f[379] && !f[329] && f[331] && !f[604];
	assign leaf[2332] = f[379] && !f[329] && f[331] && f[604];
	assign leaf[2333] = f[379] && f[329] && !f[268] && !f[431];
	assign leaf[2334] = f[379] && f[329] && !f[268] && f[431];
	assign leaf[2335] = f[379] && f[329] && f[268] && !f[540];
	assign leaf[2336] = f[379] && f[329] && f[268] && f[540];
	
	// Tree 151, Classifier 1, Iteration: 15
	assign leaf[2337] = !f[430] && !f[434] && !f[100] && !f[189];
	assign leaf[2338] = !f[430] && !f[434] && !f[100] && f[189];
	assign leaf[2339] = !f[430] && !f[434] && f[100] && !f[350];
	assign leaf[2340] = !f[430] && !f[434] && f[100] && f[350];
	assign leaf[2341] = !f[430] && f[434] && !f[298] && !f[486];
	assign leaf[2342] = !f[430] && f[434] && !f[298] && f[486];
	assign leaf[2343] = !f[430] && f[434] && f[298] && !f[237];
	assign leaf[2344] = !f[430] && f[434] && f[298] && f[237];
	assign leaf[2345] = f[430] && !f[349] && !f[649] && !f[715];
	assign leaf[2346] = f[430] && !f[349] && !f[649] && f[715];
	assign leaf[2347] = f[430] && !f[349] && f[649];
	assign leaf[2348] = f[430] && f[349] && !f[408] && !f[519];
	assign leaf[2349] = f[430] && f[349] && !f[408] && f[519];
	assign leaf[2350] = f[430] && f[349] && f[408] && !f[410];
	assign leaf[2351] = f[430] && f[349] && f[408] && f[410];
	
	// Tree 152, Classifier 2, Iteration: 15
	assign leaf[2352] = !f[345] && !f[348] && !f[342] && !f[455];
	assign leaf[2353] = !f[345] && !f[348] && !f[342] && f[455];
	assign leaf[2354] = !f[345] && !f[348] && f[342] && !f[398];
	assign leaf[2355] = !f[345] && !f[348] && f[342] && f[398];
	assign leaf[2356] = !f[345] && f[348] && !f[444] && !f[580];
	assign leaf[2357] = !f[345] && f[348] && !f[444] && f[580];
	assign leaf[2358] = !f[345] && f[348] && f[444] && !f[386];
	assign leaf[2359] = !f[345] && f[348] && f[444] && f[386];
	assign leaf[2360] = f[345] && !f[401] && !f[515] && !f[351];
	assign leaf[2361] = f[345] && !f[401] && !f[515] && f[351];
	assign leaf[2362] = f[345] && !f[401] && f[515] && !f[427];
	assign leaf[2363] = f[345] && !f[401] && f[515] && f[427];
	assign leaf[2364] = f[345] && f[401] && !f[290] && !f[482];
	assign leaf[2365] = f[345] && f[401] && !f[290] && f[482];
	assign leaf[2366] = f[345] && f[401] && f[290] && !f[667];
	assign leaf[2367] = f[345] && f[401] && f[290] && f[667];
	
	// Tree 153, Classifier 3, Iteration: 15
	assign leaf[2368] = !f[429] && !f[495] && !f[469] && !f[521];
	assign leaf[2369] = !f[429] && !f[495] && !f[469] && f[521];
	assign leaf[2370] = !f[429] && !f[495] && f[469] && !f[265];
	assign leaf[2371] = !f[429] && !f[495] && f[469] && f[265];
	assign leaf[2372] = !f[429] && f[495] && !f[398] && !f[262];
	assign leaf[2373] = !f[429] && f[495] && !f[398] && f[262];
	assign leaf[2374] = !f[429] && f[495] && f[398] && !f[371];
	assign leaf[2375] = !f[429] && f[495] && f[398] && f[371];
	assign leaf[2376] = f[429] && !f[511] && !f[318] && !f[343];
	assign leaf[2377] = f[429] && !f[511] && !f[318] && f[343];
	assign leaf[2378] = f[429] && !f[511] && f[318] && !f[231];
	assign leaf[2379] = f[429] && !f[511] && f[318] && f[231];
	assign leaf[2380] = f[429] && f[511] && !f[453] && !f[456];
	assign leaf[2381] = f[429] && f[511] && !f[453] && f[456];
	assign leaf[2382] = f[429] && f[511] && f[453] && !f[464];
	assign leaf[2383] = f[429] && f[511] && f[453] && f[464];
	
	// Tree 154, Classifier 4, Iteration: 15
	assign leaf[2384] = !f[427] && !f[375] && !f[293] && !f[209];
	assign leaf[2385] = !f[427] && !f[375] && !f[293] && f[209];
	assign leaf[2386] = !f[427] && !f[375] && f[293] && !f[190];
	assign leaf[2387] = !f[427] && !f[375] && f[293] && f[190];
	assign leaf[2388] = !f[427] && f[375] && !f[408] && !f[409];
	assign leaf[2389] = !f[427] && f[375] && !f[408] && f[409];
	assign leaf[2390] = !f[427] && f[375] && f[408] && !f[601];
	assign leaf[2391] = !f[427] && f[375] && f[408] && f[601];
	assign leaf[2392] = f[427] && !f[346] && !f[237] && !f[181];
	assign leaf[2393] = f[427] && !f[346] && !f[237] && f[181];
	assign leaf[2394] = f[427] && !f[346] && f[237] && !f[191];
	assign leaf[2395] = f[427] && !f[346] && f[237] && f[191];
	assign leaf[2396] = f[427] && f[346] && !f[328] && !f[325];
	assign leaf[2397] = f[427] && f[346] && !f[328] && f[325];
	assign leaf[2398] = f[427] && f[346] && f[328] && !f[241];
	assign leaf[2399] = f[427] && f[346] && f[328] && f[241];
	
	// Tree 155, Classifier 5, Iteration: 15
	assign leaf[2400] = !f[490] && !f[235] && !f[247] && !f[261];
	assign leaf[2401] = !f[490] && !f[235] && !f[247] && f[261];
	assign leaf[2402] = !f[490] && !f[235] && f[247] && !f[387];
	assign leaf[2403] = !f[490] && !f[235] && f[247] && f[387];
	assign leaf[2404] = !f[490] && f[235] && !f[299] && !f[330];
	assign leaf[2405] = !f[490] && f[235] && !f[299] && f[330];
	assign leaf[2406] = !f[490] && f[235] && f[299] && !f[294];
	assign leaf[2407] = !f[490] && f[235] && f[299] && f[294];
	assign leaf[2408] = f[490] && !f[380] && !f[438] && !f[350];
	assign leaf[2409] = f[490] && !f[380] && !f[438] && f[350];
	assign leaf[2410] = f[490] && !f[380] && f[438] && !f[686];
	assign leaf[2411] = f[490] && !f[380] && f[438] && f[686];
	assign leaf[2412] = f[490] && f[380] && !f[538] && !f[247];
	assign leaf[2413] = f[490] && f[380] && !f[538] && f[247];
	assign leaf[2414] = f[490] && f[380] && f[538] && !f[354];
	assign leaf[2415] = f[490] && f[380] && f[538] && f[354];
	
	// Tree 156, Classifier 6, Iteration: 15
	assign leaf[2416] = !f[414] && !f[430] && !f[416] && !f[431];
	assign leaf[2417] = !f[414] && !f[430] && !f[416] && f[431];
	assign leaf[2418] = !f[414] && !f[430] && f[416] && !f[265];
	assign leaf[2419] = !f[414] && !f[430] && f[416] && f[265];
	assign leaf[2420] = !f[414] && f[430] && !f[347] && !f[210];
	assign leaf[2421] = !f[414] && f[430] && !f[347] && f[210];
	assign leaf[2422] = !f[414] && f[430] && f[347] && !f[299];
	assign leaf[2423] = !f[414] && f[430] && f[347] && f[299];
	assign leaf[2424] = f[414] && !f[657] && !f[239] && !f[187];
	assign leaf[2425] = f[414] && !f[657] && !f[239] && f[187];
	assign leaf[2426] = f[414] && !f[657] && f[239] && !f[347];
	assign leaf[2427] = f[414] && !f[657] && f[239] && f[347];
	assign leaf[2428] = f[414] && f[657] && !f[454];
	assign leaf[2429] = f[414] && f[657] && f[454] && !f[434];
	assign leaf[2430] = f[414] && f[657] && f[454] && f[434];
	
	// Tree 157, Classifier 7, Iteration: 15
	assign leaf[2431] = !f[744] && !f[578] && !f[437] && !f[711];
	assign leaf[2432] = !f[744] && !f[578] && !f[437] && f[711];
	assign leaf[2433] = !f[744] && !f[578] && f[437] && !f[296];
	assign leaf[2434] = !f[744] && !f[578] && f[437] && f[296];
	assign leaf[2435] = !f[744] && f[578] && !f[717] && !f[340];
	assign leaf[2436] = !f[744] && f[578] && !f[717] && f[340];
	assign leaf[2437] = !f[744] && f[578] && f[717] && !f[460];
	assign leaf[2438] = !f[744] && f[578] && f[717] && f[460];
	assign leaf[2439] = f[744] && !f[461] && !f[349] && !f[374];
	assign leaf[2440] = f[744] && !f[461] && !f[349] && f[374];
	assign leaf[2441] = f[744] && !f[461] && f[349] && !f[238];
	assign leaf[2442] = f[744] && !f[461] && f[349] && f[238];
	assign leaf[2443] = f[744] && f[461] && !f[458] && !f[518];
	assign leaf[2444] = f[744] && f[461] && !f[458] && f[518];
	assign leaf[2445] = f[744] && f[461] && f[458] && !f[344];
	assign leaf[2446] = f[744] && f[461] && f[458] && f[344];
	
	// Tree 158, Classifier 8, Iteration: 15
	assign leaf[2447] = !f[467] && !f[658] && !f[513] && !f[663];
	assign leaf[2448] = !f[467] && !f[658] && !f[513] && f[663];
	assign leaf[2449] = !f[467] && !f[658] && f[513] && !f[628];
	assign leaf[2450] = !f[467] && !f[658] && f[513] && f[628];
	assign leaf[2451] = !f[467] && f[658] && !f[602] && !f[572];
	assign leaf[2452] = !f[467] && f[658] && !f[602] && f[572];
	assign leaf[2453] = !f[467] && f[658] && f[602] && !f[267];
	assign leaf[2454] = !f[467] && f[658] && f[602] && f[267];
	assign leaf[2455] = f[467] && !f[521] && !f[638] && !f[261];
	assign leaf[2456] = f[467] && !f[521] && !f[638] && f[261];
	assign leaf[2457] = f[467] && !f[521] && f[638] && !f[551];
	assign leaf[2458] = f[467] && !f[521] && f[638] && f[551];
	assign leaf[2459] = f[467] && f[521] && !f[351] && !f[637];
	assign leaf[2460] = f[467] && f[521] && !f[351] && f[637];
	assign leaf[2461] = f[467] && f[521] && f[351] && !f[274];
	assign leaf[2462] = f[467] && f[521] && f[351] && f[274];
	
	// Tree 159, Classifier 9, Iteration: 15
	assign leaf[2463] = !f[128] && !f[443] && !f[189] && !f[355];
	assign leaf[2464] = !f[128] && !f[443] && !f[189] && f[355];
	assign leaf[2465] = !f[128] && !f[443] && f[189] && !f[383];
	assign leaf[2466] = !f[128] && !f[443] && f[189] && f[383];
	assign leaf[2467] = !f[128] && f[443] && !f[639] && !f[368];
	assign leaf[2468] = !f[128] && f[443] && !f[639] && f[368];
	assign leaf[2469] = !f[128] && f[443] && f[639];
	assign leaf[2470] = f[128] && !f[275] && !f[659] && !f[358];
	assign leaf[2471] = f[128] && !f[275] && !f[659] && f[358];
	assign leaf[2472] = f[128] && !f[275] && f[659] && !f[432];
	assign leaf[2473] = f[128] && !f[275] && f[659] && f[432];
	assign leaf[2474] = f[128] && f[275];
	
	// Tree 160, Classifier 0, Iteration: 16
	assign leaf[2475] = !f[482] && !f[485] && !f[486] && !f[480];
	assign leaf[2476] = !f[482] && !f[485] && !f[486] && f[480];
	assign leaf[2477] = !f[482] && !f[485] && f[486] && !f[154];
	assign leaf[2478] = !f[482] && !f[485] && f[486] && f[154];
	assign leaf[2479] = !f[482] && f[485] && !f[656] && !f[600];
	assign leaf[2480] = !f[482] && f[485] && !f[656] && f[600];
	assign leaf[2481] = !f[482] && f[485] && f[656] && !f[541];
	assign leaf[2482] = !f[482] && f[485] && f[656] && f[541];
	assign leaf[2483] = f[482] && !f[399] && !f[516] && !f[462];
	assign leaf[2484] = f[482] && !f[399] && !f[516] && f[462];
	assign leaf[2485] = f[482] && !f[399] && f[516] && !f[219];
	assign leaf[2486] = f[482] && !f[399] && f[516] && f[219];
	assign leaf[2487] = f[482] && f[399] && !f[409] && !f[691];
	assign leaf[2488] = f[482] && f[399] && !f[409] && f[691];
	assign leaf[2489] = f[482] && f[399] && f[409] && !f[320];
	assign leaf[2490] = f[482] && f[399] && f[409] && f[320];
	
	// Tree 161, Classifier 1, Iteration: 16
	assign leaf[2491] = !f[317] && !f[628] && !f[684] && !f[204];
	assign leaf[2492] = !f[317] && !f[628] && !f[684] && f[204];
	assign leaf[2493] = !f[317] && !f[628] && f[684] && !f[631];
	assign leaf[2494] = !f[317] && !f[628] && f[684] && f[631];
	assign leaf[2495] = !f[317] && f[628] && !f[545] && !f[405];
	assign leaf[2496] = !f[317] && f[628] && !f[545] && f[405];
	assign leaf[2497] = !f[317] && f[628] && f[545] && !f[295];
	assign leaf[2498] = !f[317] && f[628] && f[545] && f[295];
	assign leaf[2499] = f[317] && !f[98] && !f[99] && !f[131];
	assign leaf[2500] = f[317] && !f[98] && !f[99] && f[131];
	assign leaf[2501] = f[317] && !f[98] && f[99];
	assign leaf[2502] = f[317] && f[98] && !f[237];
	assign leaf[2503] = f[317] && f[98] && f[237];
	
	// Tree 162, Classifier 2, Iteration: 16
	assign leaf[2504] = !f[150] && !f[657] && !f[157] && !f[471];
	assign leaf[2505] = !f[150] && !f[657] && !f[157] && f[471];
	assign leaf[2506] = !f[150] && !f[657] && f[157] && !f[322];
	assign leaf[2507] = !f[150] && !f[657] && f[157] && f[322];
	assign leaf[2508] = !f[150] && f[657] && !f[403] && !f[663];
	assign leaf[2509] = !f[150] && f[657] && !f[403] && f[663];
	assign leaf[2510] = !f[150] && f[657] && f[403] && !f[125];
	assign leaf[2511] = !f[150] && f[657] && f[403] && f[125];
	assign leaf[2512] = f[150] && !f[290] && !f[315] && !f[409];
	assign leaf[2513] = f[150] && !f[290] && !f[315] && f[409];
	assign leaf[2514] = f[150] && !f[290] && f[315] && !f[399];
	assign leaf[2515] = f[150] && !f[290] && f[315] && f[399];
	assign leaf[2516] = f[150] && f[290] && !f[269] && !f[538];
	assign leaf[2517] = f[150] && f[290] && !f[269] && f[538];
	assign leaf[2518] = f[150] && f[290] && f[269] && !f[625];
	assign leaf[2519] = f[150] && f[290] && f[269] && f[625];
	
	// Tree 163, Classifier 3, Iteration: 16
	assign leaf[2520] = !f[372] && !f[212] && !f[173] && !f[487];
	assign leaf[2521] = !f[372] && !f[212] && !f[173] && f[487];
	assign leaf[2522] = !f[372] && !f[212] && f[173] && !f[493];
	assign leaf[2523] = !f[372] && !f[212] && f[173] && f[493];
	assign leaf[2524] = !f[372] && f[212] && !f[319] && !f[405];
	assign leaf[2525] = !f[372] && f[212] && !f[319] && f[405];
	assign leaf[2526] = !f[372] && f[212] && f[319] && !f[294];
	assign leaf[2527] = !f[372] && f[212] && f[319] && f[294];
	assign leaf[2528] = f[372] && !f[321] && !f[492] && !f[259];
	assign leaf[2529] = f[372] && !f[321] && !f[492] && f[259];
	assign leaf[2530] = f[372] && !f[321] && f[492] && !f[650];
	assign leaf[2531] = f[372] && !f[321] && f[492] && f[650];
	assign leaf[2532] = f[372] && f[321] && !f[455] && !f[288];
	assign leaf[2533] = f[372] && f[321] && !f[455] && f[288];
	assign leaf[2534] = f[372] && f[321] && f[455] && !f[202];
	assign leaf[2535] = f[372] && f[321] && f[455] && f[202];
	
	// Tree 164, Classifier 4, Iteration: 16
	assign leaf[2536] = !f[568] && !f[454] && !f[375] && !f[401];
	assign leaf[2537] = !f[568] && !f[454] && !f[375] && f[401];
	assign leaf[2538] = !f[568] && !f[454] && f[375] && !f[551];
	assign leaf[2539] = !f[568] && !f[454] && f[375] && f[551];
	assign leaf[2540] = !f[568] && f[454] && !f[331] && !f[345];
	assign leaf[2541] = !f[568] && f[454] && !f[331] && f[345];
	assign leaf[2542] = !f[568] && f[454] && f[331] && !f[209];
	assign leaf[2543] = !f[568] && f[454] && f[331] && f[209];
	assign leaf[2544] = f[568] && !f[626] && !f[636] && !f[298];
	assign leaf[2545] = f[568] && !f[626] && !f[636] && f[298];
	assign leaf[2546] = f[568] && !f[626] && f[636] && !f[182];
	assign leaf[2547] = f[568] && !f[626] && f[636] && f[182];
	assign leaf[2548] = f[568] && f[626] && !f[399];
	assign leaf[2549] = f[568] && f[626] && f[399] && !f[628];
	assign leaf[2550] = f[568] && f[626] && f[399] && f[628];
	
	// Tree 165, Classifier 5, Iteration: 16
	assign leaf[2551] = !f[435] && !f[493] && !f[289] && !f[379];
	assign leaf[2552] = !f[435] && !f[493] && !f[289] && f[379];
	assign leaf[2553] = !f[435] && !f[493] && f[289] && !f[387];
	assign leaf[2554] = !f[435] && !f[493] && f[289] && f[387];
	assign leaf[2555] = !f[435] && f[493] && !f[328] && !f[216];
	assign leaf[2556] = !f[435] && f[493] && !f[328] && f[216];
	assign leaf[2557] = !f[435] && f[493] && f[328] && !f[133];
	assign leaf[2558] = !f[435] && f[493] && f[328] && f[133];
	assign leaf[2559] = f[435] && !f[353] && !f[383] && !f[323];
	assign leaf[2560] = f[435] && !f[353] && !f[383] && f[323];
	assign leaf[2561] = f[435] && !f[353] && f[383] && !f[468];
	assign leaf[2562] = f[435] && !f[353] && f[383] && f[468];
	assign leaf[2563] = f[435] && f[353] && !f[333] && !f[191];
	assign leaf[2564] = f[435] && f[353] && !f[333] && f[191];
	assign leaf[2565] = f[435] && f[353] && f[333];
	
	// Tree 166, Classifier 6, Iteration: 16
	assign leaf[2566] = !f[685] && !f[574] && !f[131] && !f[268];
	assign leaf[2567] = !f[685] && !f[574] && !f[131] && f[268];
	assign leaf[2568] = !f[685] && !f[574] && f[131] && !f[265];
	assign leaf[2569] = !f[685] && !f[574] && f[131] && f[265];
	assign leaf[2570] = !f[685] && f[574] && !f[210] && !f[156];
	assign leaf[2571] = !f[685] && f[574] && !f[210] && f[156];
	assign leaf[2572] = !f[685] && f[574] && f[210] && !f[100];
	assign leaf[2573] = !f[685] && f[574] && f[210] && f[100];
	assign leaf[2574] = f[685] && !f[192];
	assign leaf[2575] = f[685] && f[192];
	
	// Tree 167, Classifier 7, Iteration: 16
	assign leaf[2576] = !f[376] && !f[607] && !f[402] && !f[427];
	assign leaf[2577] = !f[376] && !f[607] && !f[402] && f[427];
	assign leaf[2578] = !f[376] && !f[607] && f[402] && !f[431];
	assign leaf[2579] = !f[376] && !f[607] && f[402] && f[431];
	assign leaf[2580] = !f[376] && f[607] && !f[435] && !f[717];
	assign leaf[2581] = !f[376] && f[607] && !f[435] && f[717];
	assign leaf[2582] = !f[376] && f[607] && f[435] && !f[227];
	assign leaf[2583] = !f[376] && f[607] && f[435] && f[227];
	assign leaf[2584] = f[376] && !f[384] && !f[410] && !f[740];
	assign leaf[2585] = f[376] && !f[384] && !f[410] && f[740];
	assign leaf[2586] = f[376] && !f[384] && f[410] && !f[349];
	assign leaf[2587] = f[376] && !f[384] && f[410] && f[349];
	assign leaf[2588] = f[376] && f[384] && !f[183] && !f[569];
	assign leaf[2589] = f[376] && f[384] && !f[183] && f[569];
	assign leaf[2590] = f[376] && f[384] && f[183] && !f[715];
	assign leaf[2591] = f[376] && f[384] && f[183] && f[715];
	
	// Tree 168, Classifier 8, Iteration: 16
	assign leaf[2592] = !f[434] && !f[520] && !f[549] && !f[457];
	assign leaf[2593] = !f[434] && !f[520] && !f[549] && f[457];
	assign leaf[2594] = !f[434] && !f[520] && f[549] && !f[407];
	assign leaf[2595] = !f[434] && !f[520] && f[549] && f[407];
	assign leaf[2596] = !f[434] && f[520] && !f[378] && !f[304];
	assign leaf[2597] = !f[434] && f[520] && !f[378] && f[304];
	assign leaf[2598] = !f[434] && f[520] && f[378] && !f[346];
	assign leaf[2599] = !f[434] && f[520] && f[378] && f[346];
	assign leaf[2600] = f[434] && !f[437] && !f[124] && !f[496];
	assign leaf[2601] = f[434] && !f[437] && !f[124] && f[496];
	assign leaf[2602] = f[434] && !f[437] && f[124] && !f[465];
	assign leaf[2603] = f[434] && !f[437] && f[124] && f[465];
	assign leaf[2604] = f[434] && f[437] && !f[634] && !f[541];
	assign leaf[2605] = f[434] && f[437] && !f[634] && f[541];
	assign leaf[2606] = f[434] && f[437] && f[634] && !f[315];
	assign leaf[2607] = f[434] && f[437] && f[634] && f[315];
	
	// Tree 169, Classifier 9, Iteration: 16
	assign leaf[2608] = !f[160] && !f[176] && !f[126] && !f[219];
	assign leaf[2609] = !f[160] && !f[176] && !f[126] && f[219];
	assign leaf[2610] = !f[160] && !f[176] && f[126] && !f[462];
	assign leaf[2611] = !f[160] && !f[176] && f[126] && f[462];
	assign leaf[2612] = !f[160] && f[176] && !f[694] && !f[342];
	assign leaf[2613] = !f[160] && f[176] && !f[694] && f[342];
	assign leaf[2614] = !f[160] && f[176] && f[694] && !f[440];
	assign leaf[2615] = !f[160] && f[176] && f[694] && f[440];
	assign leaf[2616] = f[160] && !f[427] && !f[572] && !f[509];
	assign leaf[2617] = f[160] && !f[427] && !f[572] && f[509];
	assign leaf[2618] = f[160] && !f[427] && f[572] && !f[318];
	assign leaf[2619] = f[160] && !f[427] && f[572] && f[318];
	assign leaf[2620] = f[160] && f[427] && !f[264];
	assign leaf[2621] = f[160] && f[427] && f[264] && !f[595];
	assign leaf[2622] = f[160] && f[427] && f[264] && f[595];
	
	// Tree 170, Classifier 0, Iteration: 17
	assign leaf[2623] = !f[406] && !f[387] && !f[402] && !f[400];
	assign leaf[2624] = !f[406] && !f[387] && !f[402] && f[400];
	assign leaf[2625] = !f[406] && !f[387] && f[402] && !f[299];
	assign leaf[2626] = !f[406] && !f[387] && f[402] && f[299];
	assign leaf[2627] = !f[406] && f[387] && !f[510] && !f[398];
	assign leaf[2628] = !f[406] && f[387] && !f[510] && f[398];
	assign leaf[2629] = !f[406] && f[387] && f[510] && !f[437];
	assign leaf[2630] = !f[406] && f[387] && f[510] && f[437];
	assign leaf[2631] = f[406] && !f[244] && !f[405] && !f[356];
	assign leaf[2632] = f[406] && !f[244] && !f[405] && f[356];
	assign leaf[2633] = f[406] && !f[244] && f[405] && !f[621];
	assign leaf[2634] = f[406] && !f[244] && f[405] && f[621];
	assign leaf[2635] = f[406] && f[244] && !f[540] && !f[508];
	assign leaf[2636] = f[406] && f[244] && !f[540] && f[508];
	assign leaf[2637] = f[406] && f[244] && f[540] && !f[357];
	assign leaf[2638] = f[406] && f[244] && f[540] && f[357];
	
	// Tree 171, Classifier 1, Iteration: 17
	assign leaf[2639] = !f[374] && !f[456] && !f[685] && !f[628];
	assign leaf[2640] = !f[374] && !f[456] && !f[685] && f[628];
	assign leaf[2641] = !f[374] && !f[456] && f[685] && !f[208];
	assign leaf[2642] = !f[374] && !f[456] && f[685] && f[208];
	assign leaf[2643] = !f[374] && f[456] && !f[376];
	assign leaf[2644] = !f[374] && f[456] && f[376] && !f[572];
	assign leaf[2645] = !f[374] && f[456] && f[376] && f[572];
	assign leaf[2646] = f[374] && !f[294];
	assign leaf[2647] = f[374] && f[294] && !f[126] && !f[687];
	assign leaf[2648] = f[374] && f[294] && !f[126] && f[687];
	assign leaf[2649] = f[374] && f[294] && f[126] && !f[491];
	assign leaf[2650] = f[374] && f[294] && f[126] && f[491];
	
	// Tree 172, Classifier 2, Iteration: 17
	assign leaf[2651] = !f[514] && !f[379] && !f[319] && !f[546];
	assign leaf[2652] = !f[514] && !f[379] && !f[319] && f[546];
	assign leaf[2653] = !f[514] && !f[379] && f[319] && !f[570];
	assign leaf[2654] = !f[514] && !f[379] && f[319] && f[570];
	assign leaf[2655] = !f[514] && f[379] && !f[516] && !f[454];
	assign leaf[2656] = !f[514] && f[379] && !f[516] && f[454];
	assign leaf[2657] = !f[514] && f[379] && f[516] && !f[607];
	assign leaf[2658] = !f[514] && f[379] && f[516] && f[607];
	assign leaf[2659] = f[514] && !f[343] && !f[580] && !f[635];
	assign leaf[2660] = f[514] && !f[343] && !f[580] && f[635];
	assign leaf[2661] = f[514] && !f[343] && f[580] && !f[468];
	assign leaf[2662] = f[514] && !f[343] && f[580] && f[468];
	assign leaf[2663] = f[514] && f[343] && !f[427] && !f[401];
	assign leaf[2664] = f[514] && f[343] && !f[427] && f[401];
	assign leaf[2665] = f[514] && f[343] && f[427] && !f[375];
	assign leaf[2666] = f[514] && f[343] && f[427] && f[375];
	
	// Tree 173, Classifier 3, Iteration: 17
	assign leaf[2667] = !f[427] && !f[202] && !f[292] && !f[317];
	assign leaf[2668] = !f[427] && !f[202] && !f[292] && f[317];
	assign leaf[2669] = !f[427] && !f[202] && f[292] && !f[267];
	assign leaf[2670] = !f[427] && !f[202] && f[292] && f[267];
	assign leaf[2671] = !f[427] && f[202] && !f[580] && !f[492];
	assign leaf[2672] = !f[427] && f[202] && !f[580] && f[492];
	assign leaf[2673] = !f[427] && f[202] && f[580] && !f[237];
	assign leaf[2674] = !f[427] && f[202] && f[580] && f[237];
	assign leaf[2675] = f[427] && !f[357] && !f[681] && !f[128];
	assign leaf[2676] = f[427] && !f[357] && !f[681] && f[128];
	assign leaf[2677] = f[427] && !f[357] && f[681] && !f[318];
	assign leaf[2678] = f[427] && !f[357] && f[681] && f[318];
	assign leaf[2679] = f[427] && f[357] && !f[189] && !f[229];
	assign leaf[2680] = f[427] && f[357] && !f[189] && f[229];
	assign leaf[2681] = f[427] && f[357] && f[189] && !f[400];
	assign leaf[2682] = f[427] && f[357] && f[189] && f[400];
	
	// Tree 174, Classifier 4, Iteration: 17
	assign leaf[2683] = !f[463] && !f[628] && !f[323] && !f[574];
	assign leaf[2684] = !f[463] && !f[628] && !f[323] && f[574];
	assign leaf[2685] = !f[463] && !f[628] && f[323] && !f[380];
	assign leaf[2686] = !f[463] && !f[628] && f[323] && f[380];
	assign leaf[2687] = !f[463] && f[628] && !f[462] && !f[219];
	assign leaf[2688] = !f[463] && f[628] && !f[462] && f[219];
	assign leaf[2689] = !f[463] && f[628] && f[462] && !f[347];
	assign leaf[2690] = !f[463] && f[628] && f[462] && f[347];
	assign leaf[2691] = f[463] && !f[740] && !f[542] && !f[208];
	assign leaf[2692] = f[463] && !f[740] && !f[542] && f[208];
	assign leaf[2693] = f[463] && !f[740] && f[542] && !f[163];
	assign leaf[2694] = f[463] && !f[740] && f[542] && f[163];
	assign leaf[2695] = f[463] && f[740] && !f[426];
	assign leaf[2696] = f[463] && f[740] && f[426];
	
	// Tree 175, Classifier 5, Iteration: 17
	assign leaf[2697] = !f[435] && !f[464] && !f[455] && !f[289];
	assign leaf[2698] = !f[435] && !f[464] && !f[455] && f[289];
	assign leaf[2699] = !f[435] && !f[464] && f[455] && !f[522];
	assign leaf[2700] = !f[435] && !f[464] && f[455] && f[522];
	assign leaf[2701] = !f[435] && f[464] && !f[383] && !f[468];
	assign leaf[2702] = !f[435] && f[464] && !f[383] && f[468];
	assign leaf[2703] = !f[435] && f[464] && f[383] && !f[509];
	assign leaf[2704] = !f[435] && f[464] && f[383] && f[509];
	assign leaf[2705] = f[435] && !f[353] && !f[383] && !f[244];
	assign leaf[2706] = f[435] && !f[353] && !f[383] && f[244];
	assign leaf[2707] = f[435] && !f[353] && f[383] && !f[497];
	assign leaf[2708] = f[435] && !f[353] && f[383] && f[497];
	assign leaf[2709] = f[435] && f[353] && !f[276] && !f[191];
	assign leaf[2710] = f[435] && f[353] && !f[276] && f[191];
	assign leaf[2711] = f[435] && f[353] && f[276] && !f[324];
	assign leaf[2712] = f[435] && f[353] && f[276] && f[324];
	
	// Tree 176, Classifier 6, Iteration: 17
	assign leaf[2713] = !f[685] && !f[623] && !f[575] && !f[269];
	assign leaf[2714] = !f[685] && !f[623] && !f[575] && f[269];
	assign leaf[2715] = !f[685] && !f[623] && f[575] && !f[631];
	assign leaf[2716] = !f[685] && !f[623] && f[575] && f[631];
	assign leaf[2717] = !f[685] && f[623] && !f[400] && !f[343];
	assign leaf[2718] = !f[685] && f[623] && !f[400] && f[343];
	assign leaf[2719] = !f[685] && f[623] && f[400] && !f[273];
	assign leaf[2720] = !f[685] && f[623] && f[400] && f[273];
	assign leaf[2721] = f[685] && !f[598];
	assign leaf[2722] = f[685] && f[598] && !f[234] && !f[158];
	assign leaf[2723] = f[685] && f[598] && !f[234] && f[158];
	assign leaf[2724] = f[685] && f[598] && f[234];
	
	// Tree 177, Classifier 7, Iteration: 17
	assign leaf[2725] = !f[159] && !f[298] && !f[348] && !f[296];
	assign leaf[2726] = !f[159] && !f[298] && !f[348] && f[296];
	assign leaf[2727] = !f[159] && !f[298] && f[348] && !f[340];
	assign leaf[2728] = !f[159] && !f[298] && f[348] && f[340];
	assign leaf[2729] = !f[159] && f[298] && !f[266] && !f[294];
	assign leaf[2730] = !f[159] && f[298] && !f[266] && f[294];
	assign leaf[2731] = !f[159] && f[298] && f[266] && !f[553];
	assign leaf[2732] = !f[159] && f[298] && f[266] && f[553];
	assign leaf[2733] = f[159] && !f[149];
	assign leaf[2734] = f[159] && f[149];
	
	// Tree 178, Classifier 8, Iteration: 17
	assign leaf[2735] = !f[440] && !f[357] && !f[410] && !f[289];
	assign leaf[2736] = !f[440] && !f[357] && !f[410] && f[289];
	assign leaf[2737] = !f[440] && !f[357] && f[410] && !f[465];
	assign leaf[2738] = !f[440] && !f[357] && f[410] && f[465];
	assign leaf[2739] = !f[440] && f[357] && !f[327] && !f[469];
	assign leaf[2740] = !f[440] && f[357] && !f[327] && f[469];
	assign leaf[2741] = !f[440] && f[357] && f[327] && !f[185];
	assign leaf[2742] = !f[440] && f[357] && f[327] && f[185];
	assign leaf[2743] = f[440] && !f[522] && !f[180] && !f[360];
	assign leaf[2744] = f[440] && !f[522] && !f[180] && f[360];
	assign leaf[2745] = f[440] && !f[522] && f[180] && !f[210];
	assign leaf[2746] = f[440] && !f[522] && f[180] && f[210];
	assign leaf[2747] = f[440] && f[522] && !f[303] && !f[611];
	assign leaf[2748] = f[440] && f[522] && !f[303] && f[611];
	assign leaf[2749] = f[440] && f[522] && f[303] && !f[399];
	assign leaf[2750] = f[440] && f[522] && f[303] && f[399];
	
	// Tree 179, Classifier 9, Iteration: 17
	assign leaf[2751] = !f[694] && !f[742] && !f[719] && !f[380];
	assign leaf[2752] = !f[694] && !f[742] && !f[719] && f[380];
	assign leaf[2753] = !f[694] && !f[742] && f[719] && !f[659];
	assign leaf[2754] = !f[694] && !f[742] && f[719] && f[659];
	assign leaf[2755] = !f[694] && f[742] && !f[259] && !f[350];
	assign leaf[2756] = !f[694] && f[742] && !f[259] && f[350];
	assign leaf[2757] = !f[694] && f[742] && f[259] && !f[329];
	assign leaf[2758] = !f[694] && f[742] && f[259] && f[329];
	assign leaf[2759] = f[694] && !f[439] && !f[465];
	assign leaf[2760] = f[694] && !f[439] && f[465] && !f[314];
	assign leaf[2761] = f[694] && !f[439] && f[465] && f[314];
	assign leaf[2762] = f[694] && f[439] && !f[174] && !f[216];
	assign leaf[2763] = f[694] && f[439] && !f[174] && f[216];
	assign leaf[2764] = f[694] && f[439] && f[174];
	
	// Tree 180, Classifier 0, Iteration: 18
	assign leaf[2765] = !f[379] && !f[518] && !f[323] && !f[462];
	assign leaf[2766] = !f[379] && !f[518] && !f[323] && f[462];
	assign leaf[2767] = !f[379] && !f[518] && f[323] && !f[238];
	assign leaf[2768] = !f[379] && !f[518] && f[323] && f[238];
	assign leaf[2769] = !f[379] && f[518] && !f[321] && !f[387];
	assign leaf[2770] = !f[379] && f[518] && !f[321] && f[387];
	assign leaf[2771] = !f[379] && f[518] && f[321] && !f[427];
	assign leaf[2772] = !f[379] && f[518] && f[321] && f[427];
	assign leaf[2773] = f[379] && !f[569] && !f[293] && !f[541];
	assign leaf[2774] = f[379] && !f[569] && !f[293] && f[541];
	assign leaf[2775] = f[379] && !f[569] && f[293] && !f[576];
	assign leaf[2776] = f[379] && !f[569] && f[293] && f[576];
	assign leaf[2777] = f[379] && f[569] && !f[377] && !f[656];
	assign leaf[2778] = f[379] && f[569] && !f[377] && f[656];
	assign leaf[2779] = f[379] && f[569] && f[377] && !f[380];
	assign leaf[2780] = f[379] && f[569] && f[377] && f[380];
	
	// Tree 181, Classifier 1, Iteration: 18
	assign leaf[2781] = !f[289] && !f[351] && !f[240] && !f[184];
	assign leaf[2782] = !f[289] && !f[351] && !f[240] && f[184];
	assign leaf[2783] = !f[289] && !f[351] && f[240] && !f[608];
	assign leaf[2784] = !f[289] && !f[351] && f[240] && f[608];
	assign leaf[2785] = !f[289] && f[351] && !f[711] && !f[510];
	assign leaf[2786] = !f[289] && f[351] && !f[711] && f[510];
	assign leaf[2787] = !f[289] && f[351] && f[711];
	assign leaf[2788] = f[289] && !f[174] && !f[98] && !f[131];
	assign leaf[2789] = f[289] && !f[174] && !f[98] && f[131];
	assign leaf[2790] = f[289] && !f[174] && f[98] && !f[293];
	assign leaf[2791] = f[289] && !f[174] && f[98] && f[293];
	assign leaf[2792] = f[289] && f[174];
	
	// Tree 182, Classifier 2, Iteration: 18
	assign leaf[2793] = !f[513] && !f[377] && !f[572] && !f[509];
	assign leaf[2794] = !f[513] && !f[377] && !f[572] && f[509];
	assign leaf[2795] = !f[513] && !f[377] && f[572] && !f[634];
	assign leaf[2796] = !f[513] && !f[377] && f[572] && f[634];
	assign leaf[2797] = !f[513] && f[377] && !f[454] && !f[487];
	assign leaf[2798] = !f[513] && f[377] && !f[454] && f[487];
	assign leaf[2799] = !f[513] && f[377] && f[454] && !f[492];
	assign leaf[2800] = !f[513] && f[377] && f[454] && f[492];
	assign leaf[2801] = f[513] && !f[370] && !f[373] && !f[348];
	assign leaf[2802] = f[513] && !f[370] && !f[373] && f[348];
	assign leaf[2803] = f[513] && !f[370] && f[373] && !f[318];
	assign leaf[2804] = f[513] && !f[370] && f[373] && f[318];
	assign leaf[2805] = f[513] && f[370] && !f[260] && !f[405];
	assign leaf[2806] = f[513] && f[370] && !f[260] && f[405];
	assign leaf[2807] = f[513] && f[370] && f[260] && !f[398];
	assign leaf[2808] = f[513] && f[370] && f[260] && f[398];
	
	// Tree 183, Classifier 3, Iteration: 18
	assign leaf[2809] = !f[551] && !f[184] && !f[581] && !f[373];
	assign leaf[2810] = !f[551] && !f[184] && !f[581] && f[373];
	assign leaf[2811] = !f[551] && !f[184] && f[581] && !f[265];
	assign leaf[2812] = !f[551] && !f[184] && f[581] && f[265];
	assign leaf[2813] = !f[551] && f[184] && !f[292] && !f[548];
	assign leaf[2814] = !f[551] && f[184] && !f[292] && f[548];
	assign leaf[2815] = !f[551] && f[184] && f[292] && !f[125];
	assign leaf[2816] = !f[551] && f[184] && f[292] && f[125];
	assign leaf[2817] = f[551] && !f[371] && !f[239] && !f[291];
	assign leaf[2818] = f[551] && !f[371] && !f[239] && f[291];
	assign leaf[2819] = f[551] && !f[371] && f[239] && !f[545];
	assign leaf[2820] = f[551] && !f[371] && f[239] && f[545];
	assign leaf[2821] = f[551] && f[371] && !f[347] && !f[400];
	assign leaf[2822] = f[551] && f[371] && !f[347] && f[400];
	assign leaf[2823] = f[551] && f[371] && f[347] && !f[482];
	assign leaf[2824] = f[551] && f[371] && f[347] && f[482];
	
	// Tree 184, Classifier 4, Iteration: 18
	assign leaf[2825] = !f[594] && !f[208] && !f[601] && !f[657];
	assign leaf[2826] = !f[594] && !f[208] && !f[601] && f[657];
	assign leaf[2827] = !f[594] && !f[208] && f[601] && !f[490];
	assign leaf[2828] = !f[594] && !f[208] && f[601] && f[490];
	assign leaf[2829] = !f[594] && f[208] && !f[184] && !f[239];
	assign leaf[2830] = !f[594] && f[208] && !f[184] && f[239];
	assign leaf[2831] = !f[594] && f[208] && f[184] && !f[183];
	assign leaf[2832] = !f[594] && f[208] && f[184] && f[183];
	assign leaf[2833] = f[594] && !f[527] && !f[372];
	assign leaf[2834] = f[594] && !f[527] && f[372] && !f[625];
	assign leaf[2835] = f[594] && !f[527] && f[372] && f[625];
	assign leaf[2836] = f[594] && f[527];
	
	// Tree 185, Classifier 5, Iteration: 18
	assign leaf[2837] = !f[277] && !f[461] && !f[130] && !f[187];
	assign leaf[2838] = !f[277] && !f[461] && !f[130] && f[187];
	assign leaf[2839] = !f[277] && !f[461] && f[130] && !f[243];
	assign leaf[2840] = !f[277] && !f[461] && f[130] && f[243];
	assign leaf[2841] = !f[277] && f[461] && !f[380] && !f[411];
	assign leaf[2842] = !f[277] && f[461] && !f[380] && f[411];
	assign leaf[2843] = !f[277] && f[461] && f[380] && !f[325];
	assign leaf[2844] = !f[277] && f[461] && f[380] && f[325];
	assign leaf[2845] = f[277] && !f[383] && !f[183] && !f[300];
	assign leaf[2846] = f[277] && !f[383] && !f[183] && f[300];
	assign leaf[2847] = f[277] && !f[383] && f[183] && !f[244];
	assign leaf[2848] = f[277] && !f[383] && f[183] && f[244];
	assign leaf[2849] = f[277] && f[383];
	
	// Tree 186, Classifier 6, Iteration: 18
	assign leaf[2850] = !f[544] && !f[570] && !f[134] && !f[119];
	assign leaf[2851] = !f[544] && !f[570] && !f[134] && f[119];
	assign leaf[2852] = !f[544] && !f[570] && f[134] && !f[241];
	assign leaf[2853] = !f[544] && !f[570] && f[134] && f[241];
	assign leaf[2854] = !f[544] && f[570] && !f[429] && !f[291];
	assign leaf[2855] = !f[544] && f[570] && !f[429] && f[291];
	assign leaf[2856] = !f[544] && f[570] && f[429] && !f[160];
	assign leaf[2857] = !f[544] && f[570] && f[429] && f[160];
	assign leaf[2858] = f[544] && !f[653] && !f[609] && !f[296];
	assign leaf[2859] = f[544] && !f[653] && !f[609] && f[296];
	assign leaf[2860] = f[544] && !f[653] && f[609] && !f[455];
	assign leaf[2861] = f[544] && !f[653] && f[609] && f[455];
	assign leaf[2862] = f[544] && f[653] && !f[132] && !f[496];
	assign leaf[2863] = f[544] && f[653] && !f[132] && f[496];
	assign leaf[2864] = f[544] && f[653] && f[132] && !f[652];
	assign leaf[2865] = f[544] && f[653] && f[132] && f[652];
	
	// Tree 187, Classifier 7, Iteration: 18
	assign leaf[2866] = !f[348] && !f[239] && !f[321] && !f[486];
	assign leaf[2867] = !f[348] && !f[239] && !f[321] && f[486];
	assign leaf[2868] = !f[348] && !f[239] && f[321] && !f[182];
	assign leaf[2869] = !f[348] && !f[239] && f[321] && f[182];
	assign leaf[2870] = !f[348] && f[239] && !f[579] && !f[234];
	assign leaf[2871] = !f[348] && f[239] && !f[579] && f[234];
	assign leaf[2872] = !f[348] && f[239] && f[579] && !f[717];
	assign leaf[2873] = !f[348] && f[239] && f[579] && f[717];
	assign leaf[2874] = f[348] && !f[328] && !f[285] && !f[266];
	assign leaf[2875] = f[348] && !f[328] && !f[285] && f[266];
	assign leaf[2876] = f[348] && !f[328] && f[285] && !f[318];
	assign leaf[2877] = f[348] && !f[328] && f[285] && f[318];
	assign leaf[2878] = f[348] && f[328] && !f[184] && !f[432];
	assign leaf[2879] = f[348] && f[328] && !f[184] && f[432];
	assign leaf[2880] = f[348] && f[328] && f[184] && !f[350];
	assign leaf[2881] = f[348] && f[328] && f[184] && f[350];
	
	// Tree 188, Classifier 8, Iteration: 18
	assign leaf[2882] = !f[434] && !f[520] && !f[457] && !f[459];
	assign leaf[2883] = !f[434] && !f[520] && !f[457] && f[459];
	assign leaf[2884] = !f[434] && !f[520] && f[457] && !f[380];
	assign leaf[2885] = !f[434] && !f[520] && f[457] && f[380];
	assign leaf[2886] = !f[434] && f[520] && !f[347] && !f[459];
	assign leaf[2887] = !f[434] && f[520] && !f[347] && f[459];
	assign leaf[2888] = !f[434] && f[520] && f[347] && !f[378];
	assign leaf[2889] = !f[434] && f[520] && f[347] && f[378];
	assign leaf[2890] = f[434] && !f[428] && !f[316] && !f[291];
	assign leaf[2891] = f[434] && !f[428] && !f[316] && f[291];
	assign leaf[2892] = f[434] && !f[428] && f[316] && !f[374];
	assign leaf[2893] = f[434] && !f[428] && f[316] && f[374];
	assign leaf[2894] = f[434] && f[428] && !f[662] && !f[595];
	assign leaf[2895] = f[434] && f[428] && !f[662] && f[595];
	assign leaf[2896] = f[434] && f[428] && f[662] && !f[573];
	assign leaf[2897] = f[434] && f[428] && f[662] && f[573];
	
	// Tree 189, Classifier 9, Iteration: 18
	assign leaf[2898] = !f[159] && !f[203] && !f[742] && !f[692];
	assign leaf[2899] = !f[159] && !f[203] && !f[742] && f[692];
	assign leaf[2900] = !f[159] && !f[203] && f[742] && !f[232];
	assign leaf[2901] = !f[159] && !f[203] && f[742] && f[232];
	assign leaf[2902] = !f[159] && f[203] && !f[314] && !f[397];
	assign leaf[2903] = !f[159] && f[203] && !f[314] && f[397];
	assign leaf[2904] = !f[159] && f[203] && f[314] && !f[206];
	assign leaf[2905] = !f[159] && f[203] && f[314] && f[206];
	assign leaf[2906] = f[159] && !f[357] && !f[346] && !f[689];
	assign leaf[2907] = f[159] && !f[357] && !f[346] && f[689];
	assign leaf[2908] = f[159] && !f[357] && f[346] && !f[549];
	assign leaf[2909] = f[159] && !f[357] && f[346] && f[549];
	assign leaf[2910] = f[159] && f[357] && !f[439];
	assign leaf[2911] = f[159] && f[357] && f[439] && !f[262];
	assign leaf[2912] = f[159] && f[357] && f[439] && f[262];
	
	// Tree 190, Classifier 0, Iteration: 19
	assign leaf[2913] = !f[570] && !f[624] && !f[543] && !f[623];
	assign leaf[2914] = !f[570] && !f[624] && !f[543] && f[623];
	assign leaf[2915] = !f[570] && !f[624] && f[543] && !f[491];
	assign leaf[2916] = !f[570] && !f[624] && f[543] && f[491];
	assign leaf[2917] = !f[570] && f[624] && !f[152] && !f[487];
	assign leaf[2918] = !f[570] && f[624] && !f[152] && f[487];
	assign leaf[2919] = !f[570] && f[624] && f[152] && !f[397];
	assign leaf[2920] = !f[570] && f[624] && f[152] && f[397];
	assign leaf[2921] = f[570] && !f[656] && !f[371] && !f[401];
	assign leaf[2922] = f[570] && !f[656] && !f[371] && f[401];
	assign leaf[2923] = f[570] && !f[656] && f[371] && !f[265];
	assign leaf[2924] = f[570] && !f[656] && f[371] && f[265];
	assign leaf[2925] = f[570] && f[656] && !f[486] && !f[456];
	assign leaf[2926] = f[570] && f[656] && !f[486] && f[456];
	assign leaf[2927] = f[570] && f[656] && f[486] && !f[608];
	assign leaf[2928] = f[570] && f[656] && f[486] && f[608];
	
	// Tree 191, Classifier 1, Iteration: 19
	assign leaf[2929] = !f[438] && !f[271] && !f[485] && !f[294];
	assign leaf[2930] = !f[438] && !f[271] && !f[485] && f[294];
	assign leaf[2931] = !f[438] && !f[271] && f[485] && !f[431];
	assign leaf[2932] = !f[438] && !f[271] && f[485] && f[431];
	assign leaf[2933] = !f[438] && f[271] && !f[183] && !f[188];
	assign leaf[2934] = !f[438] && f[271] && !f[183] && f[188];
	assign leaf[2935] = !f[438] && f[271] && f[183] && !f[409];
	assign leaf[2936] = !f[438] && f[271] && f[183] && f[409];
	assign leaf[2937] = f[438] && !f[265];
	assign leaf[2938] = f[438] && f[265] && !f[152] && !f[654];
	assign leaf[2939] = f[438] && f[265] && !f[152] && f[654];
	assign leaf[2940] = f[438] && f[265] && f[152] && !f[491];
	assign leaf[2941] = f[438] && f[265] && f[152] && f[491];
	
	// Tree 192, Classifier 2, Iteration: 19
	assign leaf[2942] = !f[373] && !f[458] && !f[377] && !f[176];
	assign leaf[2943] = !f[373] && !f[458] && !f[377] && f[176];
	assign leaf[2944] = !f[373] && !f[458] && f[377] && !f[429];
	assign leaf[2945] = !f[373] && !f[458] && f[377] && f[429];
	assign leaf[2946] = !f[373] && f[458] && !f[685] && !f[381];
	assign leaf[2947] = !f[373] && f[458] && !f[685] && f[381];
	assign leaf[2948] = !f[373] && f[458] && f[685] && !f[599];
	assign leaf[2949] = !f[373] && f[458] && f[685] && f[599];
	assign leaf[2950] = f[373] && !f[453] && !f[97] && !f[501];
	assign leaf[2951] = f[373] && !f[453] && !f[97] && f[501];
	assign leaf[2952] = f[373] && !f[453] && f[97] && !f[290];
	assign leaf[2953] = f[373] && !f[453] && f[97] && f[290];
	assign leaf[2954] = f[373] && f[453] && !f[291] && !f[295];
	assign leaf[2955] = f[373] && f[453] && !f[291] && f[295];
	assign leaf[2956] = f[373] && f[453] && f[291] && !f[581];
	assign leaf[2957] = f[373] && f[453] && f[291] && f[581];
	
	// Tree 193, Classifier 3, Iteration: 19
	assign leaf[2958] = !f[373] && !f[536] && !f[682] && !f[123];
	assign leaf[2959] = !f[373] && !f[536] && !f[682] && f[123];
	assign leaf[2960] = !f[373] && !f[536] && f[682] && !f[570];
	assign leaf[2961] = !f[373] && !f[536] && f[682] && f[570];
	assign leaf[2962] = !f[373] && f[536] && !f[327] && !f[429];
	assign leaf[2963] = !f[373] && f[536] && !f[327] && f[429];
	assign leaf[2964] = !f[373] && f[536] && f[327] && !f[458];
	assign leaf[2965] = !f[373] && f[536] && f[327] && f[458];
	assign leaf[2966] = f[373] && !f[321] && !f[345] && !f[371];
	assign leaf[2967] = f[373] && !f[321] && !f[345] && f[371];
	assign leaf[2968] = f[373] && !f[321] && f[345] && !f[200];
	assign leaf[2969] = f[373] && !f[321] && f[345] && f[200];
	assign leaf[2970] = f[373] && f[321] && !f[152] && !f[206];
	assign leaf[2971] = f[373] && f[321] && !f[152] && f[206];
	assign leaf[2972] = f[373] && f[321] && f[152] && !f[289];
	assign leaf[2973] = f[373] && f[321] && f[152] && f[289];
	
	// Tree 194, Classifier 4, Iteration: 19
	assign leaf[2974] = !f[491] && !f[629] && !f[236] && !f[180];
	assign leaf[2975] = !f[491] && !f[629] && !f[236] && f[180];
	assign leaf[2976] = !f[491] && !f[629] && f[236] && !f[291];
	assign leaf[2977] = !f[491] && !f[629] && f[236] && f[291];
	assign leaf[2978] = !f[491] && f[629] && !f[630] && !f[490];
	assign leaf[2979] = !f[491] && f[629] && !f[630] && f[490];
	assign leaf[2980] = !f[491] && f[629] && f[630] && !f[302];
	assign leaf[2981] = !f[491] && f[629] && f[630] && f[302];
	assign leaf[2982] = f[491] && !f[466] && !f[212] && !f[295];
	assign leaf[2983] = f[491] && !f[466] && !f[212] && f[295];
	assign leaf[2984] = f[491] && !f[466] && f[212] && !f[296];
	assign leaf[2985] = f[491] && !f[466] && f[212] && f[296];
	assign leaf[2986] = f[491] && f[466] && !f[260] && !f[383];
	assign leaf[2987] = f[491] && f[466] && !f[260] && f[383];
	assign leaf[2988] = f[491] && f[466] && f[260] && !f[293];
	assign leaf[2989] = f[491] && f[466] && f[260] && f[293];
	
	// Tree 195, Classifier 5, Iteration: 19
	assign leaf[2990] = !f[374] && !f[321] && !f[325] && !f[402];
	assign leaf[2991] = !f[374] && !f[321] && !f[325] && f[402];
	assign leaf[2992] = !f[374] && !f[321] && f[325] && !f[380];
	assign leaf[2993] = !f[374] && !f[321] && f[325] && f[380];
	assign leaf[2994] = !f[374] && f[321] && !f[568] && !f[187];
	assign leaf[2995] = !f[374] && f[321] && !f[568] && f[187];
	assign leaf[2996] = !f[374] && f[321] && f[568] && !f[458];
	assign leaf[2997] = !f[374] && f[321] && f[568] && f[458];
	assign leaf[2998] = f[374] && !f[456] && !f[380] && !f[410];
	assign leaf[2999] = f[374] && !f[456] && !f[380] && f[410];
	assign leaf[3000] = f[374] && !f[456] && f[380] && !f[463];
	assign leaf[3001] = f[374] && !f[456] && f[380] && f[463];
	assign leaf[3002] = f[374] && f[456] && !f[540] && !f[686];
	assign leaf[3003] = f[374] && f[456] && !f[540] && f[686];
	assign leaf[3004] = f[374] && f[456] && f[540] && !f[163];
	assign leaf[3005] = f[374] && f[456] && f[540] && f[163];
	
	// Tree 196, Classifier 6, Iteration: 19
	assign leaf[3006] = !f[522] && !f[578] && !f[132] && !f[129];
	assign leaf[3007] = !f[522] && !f[578] && !f[132] && f[129];
	assign leaf[3008] = !f[522] && !f[578] && f[132] && !f[403];
	assign leaf[3009] = !f[522] && !f[578] && f[132] && f[403];
	assign leaf[3010] = !f[522] && f[578] && !f[211] && !f[400];
	assign leaf[3011] = !f[522] && f[578] && !f[211] && f[400];
	assign leaf[3012] = !f[522] && f[578] && f[211] && !f[234];
	assign leaf[3013] = !f[522] && f[578] && f[211] && f[234];
	assign leaf[3014] = f[522] && !f[207] && !f[125] && !f[622];
	assign leaf[3015] = f[522] && !f[207] && !f[125] && f[622];
	assign leaf[3016] = f[522] && !f[207] && f[125] && !f[236];
	assign leaf[3017] = f[522] && !f[207] && f[125] && f[236];
	assign leaf[3018] = f[522] && f[207] && !f[96] && !f[414];
	assign leaf[3019] = f[522] && f[207] && !f[96] && f[414];
	assign leaf[3020] = f[522] && f[207] && f[96] && !f[183];
	assign leaf[3021] = f[522] && f[207] && f[96] && f[183];
	
	// Tree 197, Classifier 7, Iteration: 19
	assign leaf[3022] = !f[539] && !f[608] && !f[267] && !f[434];
	assign leaf[3023] = !f[539] && !f[608] && !f[267] && f[434];
	assign leaf[3024] = !f[539] && !f[608] && f[267] && !f[264];
	assign leaf[3025] = !f[539] && !f[608] && f[267] && f[264];
	assign leaf[3026] = !f[539] && f[608] && !f[746] && !f[210];
	assign leaf[3027] = !f[539] && f[608] && !f[746] && f[210];
	assign leaf[3028] = !f[539] && f[608] && f[746] && !f[207];
	assign leaf[3029] = !f[539] && f[608] && f[746] && f[207];
	assign leaf[3030] = f[539] && !f[714] && !f[229] && !f[712];
	assign leaf[3031] = f[539] && !f[714] && !f[229] && f[712];
	assign leaf[3032] = f[539] && !f[714] && f[229] && !f[569];
	assign leaf[3033] = f[539] && !f[714] && f[229] && f[569];
	assign leaf[3034] = f[539] && f[714] && !f[318];
	assign leaf[3035] = f[539] && f[714] && f[318];
	
	// Tree 198, Classifier 8, Iteration: 19
	assign leaf[3036] = !f[302] && !f[332] && !f[349] && !f[375];
	assign leaf[3037] = !f[302] && !f[332] && !f[349] && f[375];
	assign leaf[3038] = !f[302] && !f[332] && f[349] && !f[375];
	assign leaf[3039] = !f[302] && !f[332] && f[349] && f[375];
	assign leaf[3040] = !f[302] && f[332] && !f[385];
	assign leaf[3041] = !f[302] && f[332] && f[385] && !f[653];
	assign leaf[3042] = !f[302] && f[332] && f[385] && f[653];
	assign leaf[3043] = f[302] && !f[272] && !f[399] && !f[601];
	assign leaf[3044] = f[302] && !f[272] && !f[399] && f[601];
	assign leaf[3045] = f[302] && !f[272] && f[399] && !f[687];
	assign leaf[3046] = f[302] && !f[272] && f[399] && f[687];
	assign leaf[3047] = f[302] && f[272] && !f[458] && !f[296];
	assign leaf[3048] = f[302] && f[272] && !f[458] && f[296];
	assign leaf[3049] = f[302] && f[272] && f[458] && !f[352];
	assign leaf[3050] = f[302] && f[272] && f[458] && f[352];
	
	// Tree 199, Classifier 9, Iteration: 19
	assign leaf[3051] = !f[567] && !f[659] && !f[212] && !f[545];
	assign leaf[3052] = !f[567] && !f[659] && !f[212] && f[545];
	assign leaf[3053] = !f[567] && !f[659] && f[212] && !f[327];
	assign leaf[3054] = !f[567] && !f[659] && f[212] && f[327];
	assign leaf[3055] = !f[567] && f[659] && !f[545] && !f[742];
	assign leaf[3056] = !f[567] && f[659] && !f[545] && f[742];
	assign leaf[3057] = !f[567] && f[659] && f[545] && !f[485];
	assign leaf[3058] = !f[567] && f[659] && f[545] && f[485];
	assign leaf[3059] = f[567] && !f[369] && !f[485] && !f[566];
	assign leaf[3060] = f[567] && !f[369] && !f[485] && f[566];
	assign leaf[3061] = f[567] && !f[369] && f[485] && !f[399];
	assign leaf[3062] = f[567] && !f[369] && f[485] && f[399];
	assign leaf[3063] = f[567] && f[369] && !f[471] && !f[466];
	assign leaf[3064] = f[567] && f[369] && !f[471] && f[466];
	assign leaf[3065] = f[567] && f[369] && f[471];
	
	// Tree 200, Classifier 0, Iteration: 20
	assign leaf[3066] = !f[415] && !f[401] && !f[403] && !f[399];
	assign leaf[3067] = !f[415] && !f[401] && !f[403] && f[399];
	assign leaf[3068] = !f[415] && !f[401] && f[403] && !f[514];
	assign leaf[3069] = !f[415] && !f[401] && f[403] && f[514];
	assign leaf[3070] = !f[415] && f[401] && !f[484] && !f[542];
	assign leaf[3071] = !f[415] && f[401] && !f[484] && f[542];
	assign leaf[3072] = !f[415] && f[401] && f[484] && !f[654];
	assign leaf[3073] = !f[415] && f[401] && f[484] && f[654];
	assign leaf[3074] = f[415] && !f[425] && !f[275] && !f[302];
	assign leaf[3075] = f[415] && !f[425] && !f[275] && f[302];
	assign leaf[3076] = f[415] && !f[425] && f[275] && !f[319];
	assign leaf[3077] = f[415] && !f[425] && f[275] && f[319];
	assign leaf[3078] = f[415] && f[425] && !f[404] && !f[148];
	assign leaf[3079] = f[415] && f[425] && !f[404] && f[148];
	assign leaf[3080] = f[415] && f[425] && f[404] && !f[346];
	assign leaf[3081] = f[415] && f[425] && f[404] && f[346];
	
	// Tree 201, Classifier 1, Iteration: 20
	assign leaf[3082] = !f[439] && !f[683] && !f[204] && !f[537];
	assign leaf[3083] = !f[439] && !f[683] && !f[204] && f[537];
	assign leaf[3084] = !f[439] && !f[683] && f[204] && !f[625];
	assign leaf[3085] = !f[439] && !f[683] && f[204] && f[625];
	assign leaf[3086] = !f[439] && f[683] && !f[544] && !f[405];
	assign leaf[3087] = !f[439] && f[683] && !f[544] && f[405];
	assign leaf[3088] = !f[439] && f[683] && f[544] && !f[264];
	assign leaf[3089] = !f[439] && f[683] && f[544] && f[264];
	assign leaf[3090] = f[439];
	
	// Tree 202, Classifier 2, Iteration: 20
	assign leaf[3091] = !f[682] && !f[488] && !f[380] && !f[547];
	assign leaf[3092] = !f[682] && !f[488] && !f[380] && f[547];
	assign leaf[3093] = !f[682] && !f[488] && f[380] && !f[517];
	assign leaf[3094] = !f[682] && !f[488] && f[380] && f[517];
	assign leaf[3095] = !f[682] && f[488] && !f[389] && !f[508];
	assign leaf[3096] = !f[682] && f[488] && !f[389] && f[508];
	assign leaf[3097] = !f[682] && f[488] && f[389] && !f[269];
	assign leaf[3098] = !f[682] && f[488] && f[389] && f[269];
	assign leaf[3099] = f[682] && !f[658] && !f[577] && !f[387];
	assign leaf[3100] = f[682] && !f[658] && !f[577] && f[387];
	assign leaf[3101] = f[682] && !f[658] && f[577] && !f[545];
	assign leaf[3102] = f[682] && !f[658] && f[577] && f[545];
	assign leaf[3103] = f[682] && f[658] && !f[404] && !f[570];
	assign leaf[3104] = f[682] && f[658] && !f[404] && f[570];
	assign leaf[3105] = f[682] && f[658] && f[404] && !f[541];
	assign leaf[3106] = f[682] && f[658] && f[404] && f[541];
	
	// Tree 203, Classifier 3, Iteration: 20
	assign leaf[3107] = !f[578] && !f[457] && !f[625] && !f[679];
	assign leaf[3108] = !f[578] && !f[457] && !f[625] && f[679];
	assign leaf[3109] = !f[578] && !f[457] && f[625] && !f[487];
	assign leaf[3110] = !f[578] && !f[457] && f[625] && f[487];
	assign leaf[3111] = !f[578] && f[457] && !f[678] && !f[708];
	assign leaf[3112] = !f[578] && f[457] && !f[678] && f[708];
	assign leaf[3113] = !f[578] && f[457] && f[678] && !f[511];
	assign leaf[3114] = !f[578] && f[457] && f[678] && f[511];
	assign leaf[3115] = f[578] && !f[712] && !f[176] && !f[651];
	assign leaf[3116] = f[578] && !f[712] && !f[176] && f[651];
	assign leaf[3117] = f[578] && !f[712] && f[176] && !f[314];
	assign leaf[3118] = f[578] && !f[712] && f[176] && f[314];
	assign leaf[3119] = f[578] && f[712] && !f[461] && !f[372];
	assign leaf[3120] = f[578] && f[712] && !f[461] && f[372];
	assign leaf[3121] = f[578] && f[712] && f[461] && !f[206];
	assign leaf[3122] = f[578] && f[712] && f[461] && f[206];
	
	// Tree 204, Classifier 4, Iteration: 20
	assign leaf[3123] = !f[409] && !f[405] && !f[488] && !f[460];
	assign leaf[3124] = !f[409] && !f[405] && !f[488] && f[460];
	assign leaf[3125] = !f[409] && !f[405] && f[488] && !f[490];
	assign leaf[3126] = !f[409] && !f[405] && f[488] && f[490];
	assign leaf[3127] = !f[409] && f[405] && !f[521] && !f[346];
	assign leaf[3128] = !f[409] && f[405] && !f[521] && f[346];
	assign leaf[3129] = !f[409] && f[405] && f[521] && !f[410];
	assign leaf[3130] = !f[409] && f[405] && f[521] && f[410];
	assign leaf[3131] = f[409] && !f[375] && !f[265] && !f[182];
	assign leaf[3132] = f[409] && !f[375] && !f[265] && f[182];
	assign leaf[3133] = f[409] && !f[375] && f[265] && !f[426];
	assign leaf[3134] = f[409] && !f[375] && f[265] && f[426];
	assign leaf[3135] = f[409] && f[375] && !f[213] && !f[296];
	assign leaf[3136] = f[409] && f[375] && !f[213] && f[296];
	assign leaf[3137] = f[409] && f[375] && f[213] && !f[296];
	assign leaf[3138] = f[409] && f[375] && f[213] && f[296];
	
	// Tree 205, Classifier 5, Iteration: 20
	assign leaf[3139] = !f[374] && !f[292] && !f[356] && !f[325];
	assign leaf[3140] = !f[374] && !f[292] && !f[356] && f[325];
	assign leaf[3141] = !f[374] && !f[292] && f[356] && !f[471];
	assign leaf[3142] = !f[374] && !f[292] && f[356] && f[471];
	assign leaf[3143] = !f[374] && f[292] && !f[130] && !f[187];
	assign leaf[3144] = !f[374] && f[292] && !f[130] && f[187];
	assign leaf[3145] = !f[374] && f[292] && f[130] && !f[459];
	assign leaf[3146] = !f[374] && f[292] && f[130] && f[459];
	assign leaf[3147] = f[374] && !f[456] && !f[567] && !f[289];
	assign leaf[3148] = f[374] && !f[456] && !f[567] && f[289];
	assign leaf[3149] = f[374] && !f[456] && f[567] && !f[125];
	assign leaf[3150] = f[374] && !f[456] && f[567] && f[125];
	assign leaf[3151] = f[374] && f[456] && !f[686] && !f[305];
	assign leaf[3152] = f[374] && f[456] && !f[686] && f[305];
	assign leaf[3153] = f[374] && f[456] && f[686] && !f[317];
	assign leaf[3154] = f[374] && f[456] && f[686] && f[317];
	
	// Tree 206, Classifier 6, Iteration: 20
	assign leaf[3155] = !f[486] && !f[387] && !f[488] && !f[456];
	assign leaf[3156] = !f[486] && !f[387] && !f[488] && f[456];
	assign leaf[3157] = !f[486] && !f[387] && f[488] && !f[522];
	assign leaf[3158] = !f[486] && !f[387] && f[488] && f[522];
	assign leaf[3159] = !f[486] && f[387] && !f[236] && !f[291];
	assign leaf[3160] = !f[486] && f[387] && !f[236] && f[291];
	assign leaf[3161] = !f[486] && f[387] && f[236] && !f[356];
	assign leaf[3162] = !f[486] && f[387] && f[236] && f[356];
	assign leaf[3163] = f[486] && !f[430] && !f[428] && !f[485];
	assign leaf[3164] = f[486] && !f[430] && !f[428] && f[485];
	assign leaf[3165] = f[486] && !f[430] && f[428] && !f[212];
	assign leaf[3166] = f[486] && !f[430] && f[428] && f[212];
	assign leaf[3167] = f[486] && f[430] && !f[601] && !f[546];
	assign leaf[3168] = f[486] && f[430] && !f[601] && f[546];
	assign leaf[3169] = f[486] && f[430] && f[601] && !f[326];
	assign leaf[3170] = f[486] && f[430] && f[601] && f[326];
	
	// Tree 207, Classifier 7, Iteration: 20
	assign leaf[3171] = !f[376] && !f[461] && !f[515] && !f[406];
	assign leaf[3172] = !f[376] && !f[461] && !f[515] && f[406];
	assign leaf[3173] = !f[376] && !f[461] && f[515] && !f[484];
	assign leaf[3174] = !f[376] && !f[461] && f[515] && f[484];
	assign leaf[3175] = !f[376] && f[461] && !f[372] && !f[374];
	assign leaf[3176] = !f[376] && f[461] && !f[372] && f[374];
	assign leaf[3177] = !f[376] && f[461] && f[372] && !f[708];
	assign leaf[3178] = !f[376] && f[461] && f[372] && f[708];
	assign leaf[3179] = f[376] && !f[284] && !f[295] && !f[397];
	assign leaf[3180] = f[376] && !f[284] && !f[295] && f[397];
	assign leaf[3181] = f[376] && !f[284] && f[295] && !f[383];
	assign leaf[3182] = f[376] && !f[284] && f[295] && f[383];
	assign leaf[3183] = f[376] && f[284] && !f[553] && !f[271];
	assign leaf[3184] = f[376] && f[284] && !f[553] && f[271];
	assign leaf[3185] = f[376] && f[284] && f[553];
	
	// Tree 208, Classifier 8, Iteration: 20
	assign leaf[3186] = !f[441] && !f[314] && !f[401] && !f[318];
	assign leaf[3187] = !f[441] && !f[314] && !f[401] && f[318];
	assign leaf[3188] = !f[441] && !f[314] && f[401] && !f[437];
	assign leaf[3189] = !f[441] && !f[314] && f[401] && f[437];
	assign leaf[3190] = !f[441] && f[314] && !f[402] && !f[375];
	assign leaf[3191] = !f[441] && f[314] && !f[402] && f[375];
	assign leaf[3192] = !f[441] && f[314] && f[402] && !f[517];
	assign leaf[3193] = !f[441] && f[314] && f[402] && f[517];
	assign leaf[3194] = f[441] && !f[523] && !f[595] && !f[608];
	assign leaf[3195] = f[441] && !f[523] && !f[595] && f[608];
	assign leaf[3196] = f[441] && !f[523] && f[595] && !f[403];
	assign leaf[3197] = f[441] && !f[523] && f[595] && f[403];
	assign leaf[3198] = f[441] && f[523] && !f[593] && !f[691];
	assign leaf[3199] = f[441] && f[523] && !f[593] && f[691];
	assign leaf[3200] = f[441] && f[523] && f[593] && !f[330];
	assign leaf[3201] = f[441] && f[523] && f[593] && f[330];
	
	// Tree 209, Classifier 9, Iteration: 20
	assign leaf[3202] = !f[599] && !f[229] && !f[653] && !f[443];
	assign leaf[3203] = !f[599] && !f[229] && !f[653] && f[443];
	assign leaf[3204] = !f[599] && !f[229] && f[653] && !f[155];
	assign leaf[3205] = !f[599] && !f[229] && f[653] && f[155];
	assign leaf[3206] = !f[599] && f[229] && !f[177] && !f[205];
	assign leaf[3207] = !f[599] && f[229] && !f[177] && f[205];
	assign leaf[3208] = !f[599] && f[229] && f[177] && !f[183];
	assign leaf[3209] = !f[599] && f[229] && f[177] && f[183];
	assign leaf[3210] = f[599] && !f[709] && !f[680] && !f[543];
	assign leaf[3211] = f[599] && !f[709] && !f[680] && f[543];
	assign leaf[3212] = f[599] && !f[709] && f[680] && !f[207];
	assign leaf[3213] = f[599] && !f[709] && f[680] && f[207];
	assign leaf[3214] = f[599] && f[709] && !f[235] && !f[214];
	assign leaf[3215] = f[599] && f[709] && !f[235] && f[214];
	assign leaf[3216] = f[599] && f[709] && f[235] && !f[378];
	assign leaf[3217] = f[599] && f[709] && f[235] && f[378];
	
	// Tree 210, Classifier 0, Iteration: 21
	assign leaf[3218] = !f[240] && !f[350] && !f[518] && !f[214];
	assign leaf[3219] = !f[240] && !f[350] && !f[518] && f[214];
	assign leaf[3220] = !f[240] && !f[350] && f[518] && !f[442];
	assign leaf[3221] = !f[240] && !f[350] && f[518] && f[442];
	assign leaf[3222] = !f[240] && f[350] && !f[215] && !f[190];
	assign leaf[3223] = !f[240] && f[350] && !f[215] && f[190];
	assign leaf[3224] = !f[240] && f[350] && f[215] && !f[264];
	assign leaf[3225] = !f[240] && f[350] && f[215] && f[264];
	assign leaf[3226] = f[240] && !f[462] && !f[690] && !f[712];
	assign leaf[3227] = f[240] && !f[462] && !f[690] && f[712];
	assign leaf[3228] = f[240] && !f[462] && f[690] && !f[498];
	assign leaf[3229] = f[240] && !f[462] && f[690] && f[498];
	assign leaf[3230] = f[240] && f[462] && !f[512] && !f[480];
	assign leaf[3231] = f[240] && f[462] && !f[512] && f[480];
	assign leaf[3232] = f[240] && f[462] && f[512] && !f[401];
	assign leaf[3233] = f[240] && f[462] && f[512] && f[401];
	
	// Tree 211, Classifier 1, Iteration: 21
	assign leaf[3234] = !f[494] && !f[344] && !f[713] && !f[683];
	assign leaf[3235] = !f[494] && !f[344] && !f[713] && f[683];
	assign leaf[3236] = !f[494] && !f[344] && f[713] && !f[345];
	assign leaf[3237] = !f[494] && !f[344] && f[713] && f[345];
	assign leaf[3238] = !f[494] && f[344] && !f[128];
	assign leaf[3239] = !f[494] && f[344] && f[128] && !f[153];
	assign leaf[3240] = !f[494] && f[344] && f[128] && f[153];
	assign leaf[3241] = f[494] && !f[125] && !f[665] && !f[72];
	assign leaf[3242] = f[494] && !f[125] && !f[665] && f[72];
	assign leaf[3243] = f[494] && !f[125] && f[665];
	assign leaf[3244] = f[494] && f[125] && !f[237];
	assign leaf[3245] = f[494] && f[125] && f[237] && !f[459];
	assign leaf[3246] = f[494] && f[125] && f[237] && f[459];
	
	// Tree 212, Classifier 2, Iteration: 21
	assign leaf[3247] = !f[152] && !f[417] && !f[98] && !f[500];
	assign leaf[3248] = !f[152] && !f[417] && !f[98] && f[500];
	assign leaf[3249] = !f[152] && !f[417] && f[98] && !f[292];
	assign leaf[3250] = !f[152] && !f[417] && f[98] && f[292];
	assign leaf[3251] = !f[152] && f[417] && !f[343] && !f[240];
	assign leaf[3252] = !f[152] && f[417] && !f[343] && f[240];
	assign leaf[3253] = !f[152] && f[417] && f[343];
	assign leaf[3254] = f[152] && !f[291] && !f[315] && !f[637];
	assign leaf[3255] = f[152] && !f[291] && !f[315] && f[637];
	assign leaf[3256] = f[152] && !f[291] && f[315] && !f[655];
	assign leaf[3257] = f[152] && !f[291] && f[315] && f[655];
	assign leaf[3258] = f[152] && f[291] && !f[547] && !f[462];
	assign leaf[3259] = f[152] && f[291] && !f[547] && f[462];
	assign leaf[3260] = f[152] && f[291] && f[547] && !f[240];
	assign leaf[3261] = f[152] && f[291] && f[547] && f[240];
	
	// Tree 213, Classifier 3, Iteration: 21
	assign leaf[3262] = !f[429] && !f[537] && !f[544] && !f[240];
	assign leaf[3263] = !f[429] && !f[537] && !f[544] && f[240];
	assign leaf[3264] = !f[429] && !f[537] && f[544] && !f[489];
	assign leaf[3265] = !f[429] && !f[537] && f[544] && f[489];
	assign leaf[3266] = !f[429] && f[537] && !f[326] && !f[382];
	assign leaf[3267] = !f[429] && f[537] && !f[326] && f[382];
	assign leaf[3268] = !f[429] && f[537] && f[326] && !f[545];
	assign leaf[3269] = !f[429] && f[537] && f[326] && f[545];
	assign leaf[3270] = f[429] && !f[512] && !f[404] && !f[582];
	assign leaf[3271] = f[429] && !f[512] && !f[404] && f[582];
	assign leaf[3272] = f[429] && !f[512] && f[404] && !f[370];
	assign leaf[3273] = f[429] && !f[512] && f[404] && f[370];
	assign leaf[3274] = f[429] && f[512] && !f[425] && !f[484];
	assign leaf[3275] = f[429] && f[512] && !f[425] && f[484];
	assign leaf[3276] = f[429] && f[512] && f[425];
	
	// Tree 214, Classifier 4, Iteration: 21
	assign leaf[3277] = !f[491] && !f[629] && !f[322] && !f[657];
	assign leaf[3278] = !f[491] && !f[629] && !f[322] && f[657];
	assign leaf[3279] = !f[491] && !f[629] && f[322] && !f[289];
	assign leaf[3280] = !f[491] && !f[629] && f[322] && f[289];
	assign leaf[3281] = !f[491] && f[629] && !f[184] && !f[685];
	assign leaf[3282] = !f[491] && f[629] && !f[184] && f[685];
	assign leaf[3283] = !f[491] && f[629] && f[184];
	assign leaf[3284] = f[491] && !f[214] && !f[269] && !f[551];
	assign leaf[3285] = f[491] && !f[214] && !f[269] && f[551];
	assign leaf[3286] = f[491] && !f[214] && f[269] && !f[270];
	assign leaf[3287] = f[491] && !f[214] && f[269] && f[270];
	assign leaf[3288] = f[491] && f[214] && !f[297] && !f[468];
	assign leaf[3289] = f[491] && f[214] && !f[297] && f[468];
	assign leaf[3290] = f[491] && f[214] && f[297] && !f[183];
	assign leaf[3291] = f[491] && f[214] && f[297] && f[183];
	
	// Tree 215, Classifier 5, Iteration: 21
	assign leaf[3292] = !f[461] && !f[305] && !f[459] && !f[131];
	assign leaf[3293] = !f[461] && !f[305] && !f[459] && f[131];
	assign leaf[3294] = !f[461] && !f[305] && f[459] && !f[542];
	assign leaf[3295] = !f[461] && !f[305] && f[459] && f[542];
	assign leaf[3296] = !f[461] && f[305] && !f[300];
	assign leaf[3297] = !f[461] && f[305] && f[300] && !f[239];
	assign leaf[3298] = !f[461] && f[305] && f[300] && f[239];
	assign leaf[3299] = f[461] && !f[381] && !f[273] && !f[351];
	assign leaf[3300] = f[461] && !f[381] && !f[273] && f[351];
	assign leaf[3301] = f[461] && !f[381] && f[273] && !f[412];
	assign leaf[3302] = f[461] && !f[381] && f[273] && f[412];
	assign leaf[3303] = f[461] && f[381] && !f[551] && !f[536];
	assign leaf[3304] = f[461] && f[381] && !f[551] && f[536];
	assign leaf[3305] = f[461] && f[381] && f[551] && !f[657];
	assign leaf[3306] = f[461] && f[381] && f[551] && f[657];
	
	// Tree 216, Classifier 6, Iteration: 21
	assign leaf[3307] = !f[297] && !f[273] && !f[351] && !f[271];
	assign leaf[3308] = !f[297] && !f[273] && !f[351] && f[271];
	assign leaf[3309] = !f[297] && !f[273] && f[351] && !f[430];
	assign leaf[3310] = !f[297] && !f[273] && f[351] && f[430];
	assign leaf[3311] = !f[297] && f[273] && !f[121] && !f[328];
	assign leaf[3312] = !f[297] && f[273] && !f[121] && f[328];
	assign leaf[3313] = !f[297] && f[273] && f[121] && !f[326];
	assign leaf[3314] = !f[297] && f[273] && f[121] && f[326];
	assign leaf[3315] = f[297] && !f[329] && !f[331] && !f[384];
	assign leaf[3316] = f[297] && !f[329] && !f[331] && f[384];
	assign leaf[3317] = f[297] && !f[329] && f[331] && !f[245];
	assign leaf[3318] = f[297] && !f[329] && f[331] && f[245];
	assign leaf[3319] = f[297] && f[329] && !f[150] && !f[379];
	assign leaf[3320] = f[297] && f[329] && !f[150] && f[379];
	assign leaf[3321] = f[297] && f[329] && f[150] && !f[209];
	assign leaf[3322] = f[297] && f[329] && f[150] && f[209];
	
	// Tree 217, Classifier 7, Iteration: 21
	assign leaf[3323] = !f[566] && !f[270] && !f[324] && !f[678];
	assign leaf[3324] = !f[566] && !f[270] && !f[324] && f[678];
	assign leaf[3325] = !f[566] && !f[270] && f[324] && !f[570];
	assign leaf[3326] = !f[566] && !f[270] && f[324] && f[570];
	assign leaf[3327] = !f[566] && f[270] && !f[486] && !f[378];
	assign leaf[3328] = !f[566] && f[270] && !f[486] && f[378];
	assign leaf[3329] = !f[566] && f[270] && f[486] && !f[399];
	assign leaf[3330] = !f[566] && f[270] && f[486] && f[399];
	assign leaf[3331] = f[566] && !f[648] && !f[341] && !f[123];
	assign leaf[3332] = f[566] && !f[648] && !f[341] && f[123];
	assign leaf[3333] = f[566] && !f[648] && f[341];
	assign leaf[3334] = f[566] && f[648];
	
	// Tree 218, Classifier 8, Iteration: 21
	assign leaf[3335] = !f[153] && !f[186] && !f[158] && !f[542];
	assign leaf[3336] = !f[153] && !f[186] && !f[158] && f[542];
	assign leaf[3337] = !f[153] && !f[186] && f[158] && !f[326];
	assign leaf[3338] = !f[153] && !f[186] && f[158] && f[326];
	assign leaf[3339] = !f[153] && f[186] && !f[241] && !f[322];
	assign leaf[3340] = !f[153] && f[186] && !f[241] && f[322];
	assign leaf[3341] = !f[153] && f[186] && f[241] && !f[659];
	assign leaf[3342] = !f[153] && f[186] && f[241] && f[659];
	assign leaf[3343] = f[153] && !f[210] && !f[350] && !f[376];
	assign leaf[3344] = f[153] && !f[210] && !f[350] && f[376];
	assign leaf[3345] = f[153] && !f[210] && f[350] && !f[293];
	assign leaf[3346] = f[153] && !f[210] && f[350] && f[293];
	assign leaf[3347] = f[153] && f[210] && !f[289] && !f[343];
	assign leaf[3348] = f[153] && f[210] && !f[289] && f[343];
	assign leaf[3349] = f[153] && f[210] && f[289] && !f[264];
	assign leaf[3350] = f[153] && f[210] && f[289] && f[264];
	
	// Tree 219, Classifier 9, Iteration: 21
	assign leaf[3351] = !f[150] && !f[129] && !f[191] && !f[355];
	assign leaf[3352] = !f[150] && !f[129] && !f[191] && f[355];
	assign leaf[3353] = !f[150] && !f[129] && f[191] && !f[187];
	assign leaf[3354] = !f[150] && !f[129] && f[191] && f[187];
	assign leaf[3355] = !f[150] && f[129] && !f[126] && !f[609];
	assign leaf[3356] = !f[150] && f[129] && !f[126] && f[609];
	assign leaf[3357] = !f[150] && f[129] && f[126] && !f[289];
	assign leaf[3358] = !f[150] && f[129] && f[126] && f[289];
	assign leaf[3359] = f[150] && !f[259] && !f[685] && !f[686];
	assign leaf[3360] = f[150] && !f[259] && !f[685] && f[686];
	assign leaf[3361] = f[150] && !f[259] && f[685] && !f[411];
	assign leaf[3362] = f[150] && !f[259] && f[685] && f[411];
	assign leaf[3363] = f[150] && f[259] && !f[522] && !f[267];
	assign leaf[3364] = f[150] && f[259] && !f[522] && f[267];
	assign leaf[3365] = f[150] && f[259] && f[522] && !f[464];
	assign leaf[3366] = f[150] && f[259] && f[522] && f[464];
	
	// Tree 220, Classifier 0, Iteration: 22
	assign leaf[3367] = !f[453] && !f[429] && !f[431] && !f[427];
	assign leaf[3368] = !f[453] && !f[429] && !f[431] && f[427];
	assign leaf[3369] = !f[453] && !f[429] && f[431] && !f[241];
	assign leaf[3370] = !f[453] && !f[429] && f[431] && f[241];
	assign leaf[3371] = !f[453] && f[429] && !f[513] && !f[511];
	assign leaf[3372] = !f[453] && f[429] && !f[513] && f[511];
	assign leaf[3373] = !f[453] && f[429] && f[513] && !f[328];
	assign leaf[3374] = !f[453] && f[429] && f[513] && f[328];
	assign leaf[3375] = f[453] && !f[458] && !f[623] && !f[410];
	assign leaf[3376] = f[453] && !f[458] && !f[623] && f[410];
	assign leaf[3377] = f[453] && !f[458] && f[623] && !f[404];
	assign leaf[3378] = f[453] && !f[458] && f[623] && f[404];
	assign leaf[3379] = f[453] && f[458] && !f[346] && !f[470];
	assign leaf[3380] = f[453] && f[458] && !f[346] && f[470];
	assign leaf[3381] = f[453] && f[458] && f[346] && !f[544];
	assign leaf[3382] = f[453] && f[458] && f[346] && f[544];
	
	// Tree 221, Classifier 1, Iteration: 22
	assign leaf[3383] = !f[289] && !f[629] && !f[211] && !f[155];
	assign leaf[3384] = !f[289] && !f[629] && !f[211] && f[155];
	assign leaf[3385] = !f[289] && !f[629] && f[211] && !f[326];
	assign leaf[3386] = !f[289] && !f[629] && f[211] && f[326];
	assign leaf[3387] = !f[289] && f[629] && !f[545] && !f[433];
	assign leaf[3388] = !f[289] && f[629] && !f[545] && f[433];
	assign leaf[3389] = !f[289] && f[629] && f[545] && !f[294];
	assign leaf[3390] = !f[289] && f[629] && f[545] && f[294];
	assign leaf[3391] = f[289] && !f[578] && !f[606];
	assign leaf[3392] = f[289] && !f[578] && f[606];
	assign leaf[3393] = f[289] && f[578] && !f[491];
	assign leaf[3394] = f[289] && f[578] && f[491] && !f[206];
	assign leaf[3395] = f[289] && f[578] && f[491] && f[206];
	
	// Tree 222, Classifier 2, Iteration: 22
	assign leaf[3396] = !f[380] && !f[397] && !f[372] && !f[204];
	assign leaf[3397] = !f[380] && !f[397] && !f[372] && f[204];
	assign leaf[3398] = !f[380] && !f[397] && f[372] && !f[377];
	assign leaf[3399] = !f[380] && !f[397] && f[372] && f[377];
	assign leaf[3400] = !f[380] && f[397] && !f[405] && !f[451];
	assign leaf[3401] = !f[380] && f[397] && !f[405] && f[451];
	assign leaf[3402] = !f[380] && f[397] && f[405] && !f[159];
	assign leaf[3403] = !f[380] && f[397] && f[405] && f[159];
	assign leaf[3404] = f[380] && !f[438] && !f[634] && !f[579];
	assign leaf[3405] = f[380] && !f[438] && !f[634] && f[579];
	assign leaf[3406] = f[380] && !f[438] && f[634] && !f[493];
	assign leaf[3407] = f[380] && !f[438] && f[634] && f[493];
	assign leaf[3408] = f[380] && f[438] && !f[511] && !f[499];
	assign leaf[3409] = f[380] && f[438] && !f[511] && f[499];
	assign leaf[3410] = f[380] && f[438] && f[511] && !f[630];
	assign leaf[3411] = f[380] && f[438] && f[511] && f[630];
	
	// Tree 223, Classifier 3, Iteration: 22
	assign leaf[3412] = !f[373] && !f[320] && !f[406] && !f[323];
	assign leaf[3413] = !f[373] && !f[320] && !f[406] && f[323];
	assign leaf[3414] = !f[373] && !f[320] && f[406] && !f[353];
	assign leaf[3415] = !f[373] && !f[320] && f[406] && f[353];
	assign leaf[3416] = !f[373] && f[320] && !f[294] && !f[174];
	assign leaf[3417] = !f[373] && f[320] && !f[294] && f[174];
	assign leaf[3418] = !f[373] && f[320] && f[294] && !f[431];
	assign leaf[3419] = !f[373] && f[320] && f[294] && f[431];
	assign leaf[3420] = f[373] && !f[321] && !f[200] && !f[345];
	assign leaf[3421] = f[373] && !f[321] && !f[200] && f[345];
	assign leaf[3422] = f[373] && !f[321] && f[200] && !f[240];
	assign leaf[3423] = f[373] && !f[321] && f[200] && f[240];
	assign leaf[3424] = f[373] && f[321] && !f[327] && !f[246];
	assign leaf[3425] = f[373] && f[321] && !f[327] && f[246];
	assign leaf[3426] = f[373] && f[321] && f[327] && !f[455];
	assign leaf[3427] = f[373] && f[321] && f[327] && f[455];
	
	// Tree 224, Classifier 4, Iteration: 22
	assign leaf[3428] = !f[430] && !f[625] && !f[482] && !f[347];
	assign leaf[3429] = !f[430] && !f[625] && !f[482] && f[347];
	assign leaf[3430] = !f[430] && !f[625] && f[482] && !f[406];
	assign leaf[3431] = !f[430] && !f[625] && f[482] && f[406];
	assign leaf[3432] = !f[430] && f[625] && !f[406] && !f[458];
	assign leaf[3433] = !f[430] && f[625] && !f[406] && f[458];
	assign leaf[3434] = !f[430] && f[625] && f[406] && !f[186];
	assign leaf[3435] = !f[430] && f[625] && f[406] && f[186];
	assign leaf[3436] = f[430] && !f[552] && !f[462] && !f[629];
	assign leaf[3437] = f[430] && !f[552] && !f[462] && f[629];
	assign leaf[3438] = f[430] && !f[552] && f[462] && !f[214];
	assign leaf[3439] = f[430] && !f[552] && f[462] && f[214];
	assign leaf[3440] = f[430] && f[552] && !f[270] && !f[273];
	assign leaf[3441] = f[430] && f[552] && !f[270] && f[273];
	assign leaf[3442] = f[430] && f[552] && f[270] && !f[209];
	assign leaf[3443] = f[430] && f[552] && f[270] && f[209];
	
	// Tree 225, Classifier 5, Iteration: 22
	assign leaf[3444] = !f[627] && !f[304] && !f[216] && !f[273];
	assign leaf[3445] = !f[627] && !f[304] && !f[216] && f[273];
	assign leaf[3446] = !f[627] && !f[304] && f[216] && !f[300];
	assign leaf[3447] = !f[627] && !f[304] && f[216] && f[300];
	assign leaf[3448] = !f[627] && f[304] && !f[301] && !f[377];
	assign leaf[3449] = !f[627] && f[304] && !f[301] && f[377];
	assign leaf[3450] = !f[627] && f[304] && f[301] && !f[359];
	assign leaf[3451] = !f[627] && f[304] && f[301] && f[359];
	assign leaf[3452] = f[627] && !f[513] && !f[517] && !f[236];
	assign leaf[3453] = f[627] && !f[513] && !f[517] && f[236];
	assign leaf[3454] = f[627] && !f[513] && f[517] && !f[381];
	assign leaf[3455] = f[627] && !f[513] && f[517] && f[381];
	assign leaf[3456] = f[627] && f[513] && !f[458] && !f[602];
	assign leaf[3457] = f[627] && f[513] && !f[458] && f[602];
	assign leaf[3458] = f[627] && f[513] && f[458] && !f[177];
	assign leaf[3459] = f[627] && f[513] && f[458] && f[177];
	
	// Tree 226, Classifier 6, Iteration: 22
	assign leaf[3460] = !f[683] && !f[635] && !f[622] && !f[687];
	assign leaf[3461] = !f[683] && !f[635] && !f[622] && f[687];
	assign leaf[3462] = !f[683] && !f[635] && f[622] && !f[498];
	assign leaf[3463] = !f[683] && !f[635] && f[622] && f[498];
	assign leaf[3464] = !f[683] && f[635] && !f[345] && !f[518];
	assign leaf[3465] = !f[683] && f[635] && !f[345] && f[518];
	assign leaf[3466] = !f[683] && f[635] && f[345] && !f[245];
	assign leaf[3467] = !f[683] && f[635] && f[345] && f[245];
	assign leaf[3468] = f[683];
	
	// Tree 227, Classifier 7, Iteration: 22
	assign leaf[3469] = !f[437] && !f[431] && !f[744] && !f[707];
	assign leaf[3470] = !f[437] && !f[431] && !f[744] && f[707];
	assign leaf[3471] = !f[437] && !f[431] && f[744] && !f[350];
	assign leaf[3472] = !f[437] && !f[431] && f[744] && f[350];
	assign leaf[3473] = !f[437] && f[431] && !f[466] && !f[383];
	assign leaf[3474] = !f[437] && f[431] && !f[466] && f[383];
	assign leaf[3475] = !f[437] && f[431] && f[466] && !f[411];
	assign leaf[3476] = !f[437] && f[431] && f[466] && f[411];
	assign leaf[3477] = f[437] && !f[606] && !f[232] && !f[484];
	assign leaf[3478] = f[437] && !f[606] && !f[232] && f[484];
	assign leaf[3479] = f[437] && !f[606] && f[232] && !f[343];
	assign leaf[3480] = f[437] && !f[606] && f[232] && f[343];
	assign leaf[3481] = f[437] && f[606] && !f[717] && !f[284];
	assign leaf[3482] = f[437] && f[606] && !f[717] && f[284];
	assign leaf[3483] = f[437] && f[606] && f[717] && !f[516];
	assign leaf[3484] = f[437] && f[606] && f[717] && f[516];
	
	// Tree 228, Classifier 8, Iteration: 22
	assign leaf[3485] = !f[688] && !f[219] && !f[631] && !f[596];
	assign leaf[3486] = !f[688] && !f[219] && !f[631] && f[596];
	assign leaf[3487] = !f[688] && !f[219] && f[631] && !f[516];
	assign leaf[3488] = !f[688] && !f[219] && f[631] && f[516];
	assign leaf[3489] = !f[688] && f[219] && !f[400] && !f[508];
	assign leaf[3490] = !f[688] && f[219] && !f[400] && f[508];
	assign leaf[3491] = !f[688] && f[219] && f[400] && !f[347];
	assign leaf[3492] = !f[688] && f[219] && f[400] && f[347];
	assign leaf[3493] = f[688] && !f[573] && !f[571] && !f[569];
	assign leaf[3494] = f[688] && !f[573] && !f[571] && f[569];
	assign leaf[3495] = f[688] && !f[573] && f[571] && !f[630];
	assign leaf[3496] = f[688] && !f[573] && f[571] && f[630];
	assign leaf[3497] = f[688] && f[573] && !f[513] && !f[717];
	assign leaf[3498] = f[688] && f[573] && !f[513] && f[717];
	assign leaf[3499] = f[688] && f[573] && f[513] && !f[214];
	assign leaf[3500] = f[688] && f[573] && f[513] && f[214];
	
	// Tree 229, Classifier 9, Iteration: 22
	assign leaf[3501] = !f[469] && !f[353] && !f[405] && !f[455];
	assign leaf[3502] = !f[469] && !f[353] && !f[405] && f[455];
	assign leaf[3503] = !f[469] && !f[353] && f[405] && !f[660];
	assign leaf[3504] = !f[469] && !f[353] && f[405] && f[660];
	assign leaf[3505] = !f[469] && f[353] && !f[378] && !f[350];
	assign leaf[3506] = !f[469] && f[353] && !f[378] && f[350];
	assign leaf[3507] = !f[469] && f[353] && f[378] && !f[461];
	assign leaf[3508] = !f[469] && f[353] && f[378] && f[461];
	assign leaf[3509] = f[469] && !f[385] && !f[667] && !f[720];
	assign leaf[3510] = f[469] && !f[385] && !f[667] && f[720];
	assign leaf[3511] = f[469] && !f[385] && f[667];
	assign leaf[3512] = f[469] && f[385] && !f[313] && !f[470];
	assign leaf[3513] = f[469] && f[385] && !f[313] && f[470];
	assign leaf[3514] = f[469] && f[385] && f[313] && !f[182];
	assign leaf[3515] = f[469] && f[385] && f[313] && f[182];
	
	// Tree 230, Classifier 0, Iteration: 23
	assign leaf[3516] = !f[663] && !f[434] && !f[241] && !f[215];
	assign leaf[3517] = !f[663] && !f[434] && !f[241] && f[215];
	assign leaf[3518] = !f[663] && !f[434] && f[241] && !f[713];
	assign leaf[3519] = !f[663] && !f[434] && f[241] && f[713];
	assign leaf[3520] = !f[663] && f[434] && !f[540] && !f[481];
	assign leaf[3521] = !f[663] && f[434] && !f[540] && f[481];
	assign leaf[3522] = !f[663] && f[434] && f[540] && !f[328];
	assign leaf[3523] = !f[663] && f[434] && f[540] && f[328];
	assign leaf[3524] = f[663] && !f[526] && !f[546] && !f[572];
	assign leaf[3525] = f[663] && !f[526] && !f[546] && f[572];
	assign leaf[3526] = f[663] && !f[526] && f[546] && !f[464];
	assign leaf[3527] = f[663] && !f[526] && f[546] && f[464];
	assign leaf[3528] = f[663] && f[526] && !f[347] && !f[402];
	assign leaf[3529] = f[663] && f[526] && !f[347] && f[402];
	assign leaf[3530] = f[663] && f[526] && f[347] && !f[551];
	assign leaf[3531] = f[663] && f[526] && f[347] && f[551];
	
	// Tree 231, Classifier 1, Iteration: 23
	assign leaf[3532] = !f[300] && !f[440] && !f[715] && !f[242];
	assign leaf[3533] = !f[300] && !f[440] && !f[715] && f[242];
	assign leaf[3534] = !f[300] && !f[440] && f[715] && !f[429];
	assign leaf[3535] = !f[300] && !f[440] && f[715] && f[429];
	assign leaf[3536] = !f[300] && f[440];
	assign leaf[3537] = f[300] && !f[162] && !f[515];
	assign leaf[3538] = f[300] && !f[162] && f[515] && !f[266];
	assign leaf[3539] = f[300] && !f[162] && f[515] && f[266];
	assign leaf[3540] = f[300] && f[162] && !f[265] && !f[573];
	assign leaf[3541] = f[300] && f[162] && !f[265] && f[573];
	assign leaf[3542] = f[300] && f[162] && f[265];
	
	// Tree 232, Classifier 2, Iteration: 23
	assign leaf[3543] = !f[685] && !f[353] && !f[122] && !f[566];
	assign leaf[3544] = !f[685] && !f[353] && !f[122] && f[566];
	assign leaf[3545] = !f[685] && !f[353] && f[122] && !f[318];
	assign leaf[3546] = !f[685] && !f[353] && f[122] && f[318];
	assign leaf[3547] = !f[685] && f[353] && !f[322] && !f[356];
	assign leaf[3548] = !f[685] && f[353] && !f[322] && f[356];
	assign leaf[3549] = !f[685] && f[353] && f[322] && !f[582];
	assign leaf[3550] = !f[685] && f[353] && f[322] && f[582];
	assign leaf[3551] = f[685] && !f[665] && !f[717] && !f[376];
	assign leaf[3552] = f[685] && !f[665] && !f[717] && f[376];
	assign leaf[3553] = f[685] && !f[665] && f[717];
	assign leaf[3554] = f[685] && f[665] && !f[582] && !f[463];
	assign leaf[3555] = f[685] && f[665] && !f[582] && f[463];
	assign leaf[3556] = f[685] && f[665] && f[582];
	
	// Tree 233, Classifier 3, Iteration: 23
	assign leaf[3557] = !f[386] && !f[485] && !f[654] && !f[569];
	assign leaf[3558] = !f[386] && !f[485] && !f[654] && f[569];
	assign leaf[3559] = !f[386] && !f[485] && f[654] && !f[543];
	assign leaf[3560] = !f[386] && !f[485] && f[654] && f[543];
	assign leaf[3561] = !f[386] && f[485] && !f[480] && !f[710];
	assign leaf[3562] = !f[386] && f[485] && !f[480] && f[710];
	assign leaf[3563] = !f[386] && f[485] && f[480] && !f[570];
	assign leaf[3564] = !f[386] && f[485] && f[480] && f[570];
	assign leaf[3565] = f[386] && !f[355];
	assign leaf[3566] = f[386] && f[355] && !f[294] && !f[564];
	assign leaf[3567] = f[386] && f[355] && !f[294] && f[564];
	assign leaf[3568] = f[386] && f[355] && f[294] && !f[150];
	assign leaf[3569] = f[386] && f[355] && f[294] && f[150];
	
	// Tree 234, Classifier 4, Iteration: 23
	assign leaf[3570] = !f[465] && !f[577] && !f[212] && !f[295];
	assign leaf[3571] = !f[465] && !f[577] && !f[212] && f[295];
	assign leaf[3572] = !f[465] && !f[577] && f[212] && !f[237];
	assign leaf[3573] = !f[465] && !f[577] && f[212] && f[237];
	assign leaf[3574] = !f[465] && f[577] && !f[662] && !f[688];
	assign leaf[3575] = !f[465] && f[577] && !f[662] && f[688];
	assign leaf[3576] = !f[465] && f[577] && f[662] && !f[179];
	assign leaf[3577] = !f[465] && f[577] && f[662] && f[179];
	assign leaf[3578] = f[465] && !f[235] && !f[179] && !f[571];
	assign leaf[3579] = f[465] && !f[235] && !f[179] && f[571];
	assign leaf[3580] = f[465] && !f[235] && f[179] && !f[262];
	assign leaf[3581] = f[465] && !f[235] && f[179] && f[262];
	assign leaf[3582] = f[465] && f[235] && !f[232] && !f[184];
	assign leaf[3583] = f[465] && f[235] && !f[232] && f[184];
	assign leaf[3584] = f[465] && f[235] && f[232] && !f[219];
	assign leaf[3585] = f[465] && f[235] && f[232] && f[219];
	
	// Tree 235, Classifier 5, Iteration: 23
	assign leaf[3586] = !f[462] && !f[464] && !f[228] && !f[610];
	assign leaf[3587] = !f[462] && !f[464] && !f[228] && f[610];
	assign leaf[3588] = !f[462] && !f[464] && f[228] && !f[691];
	assign leaf[3589] = !f[462] && !f[464] && f[228] && f[691];
	assign leaf[3590] = !f[462] && f[464] && !f[353] && !f[411];
	assign leaf[3591] = !f[462] && f[464] && !f[353] && f[411];
	assign leaf[3592] = !f[462] && f[464] && f[353] && !f[132];
	assign leaf[3593] = !f[462] && f[464] && f[353] && f[132];
	assign leaf[3594] = f[462] && !f[353] && !f[383] && !f[271];
	assign leaf[3595] = f[462] && !f[353] && !f[383] && f[271];
	assign leaf[3596] = f[462] && !f[353] && f[383] && !f[660];
	assign leaf[3597] = f[462] && !f[353] && f[383] && f[660];
	assign leaf[3598] = f[462] && f[353] && !f[331] && !f[247];
	assign leaf[3599] = f[462] && f[353] && !f[331] && f[247];
	assign leaf[3600] = f[462] && f[353] && f[331] && !f[321];
	assign leaf[3601] = f[462] && f[353] && f[331] && f[321];
	
	// Tree 236, Classifier 6, Iteration: 23
	assign leaf[3602] = !f[325] && !f[301] && !f[351] && !f[299];
	assign leaf[3603] = !f[325] && !f[301] && !f[351] && f[299];
	assign leaf[3604] = !f[325] && !f[301] && f[351] && !f[431];
	assign leaf[3605] = !f[325] && !f[301] && f[351] && f[431];
	assign leaf[3606] = !f[325] && f[301] && !f[415] && !f[122];
	assign leaf[3607] = !f[325] && f[301] && !f[415] && f[122];
	assign leaf[3608] = !f[325] && f[301] && f[415] && !f[381];
	assign leaf[3609] = !f[325] && f[301] && f[415] && f[381];
	assign leaf[3610] = f[325] && !f[357] && !f[359] && !f[384];
	assign leaf[3611] = f[325] && !f[357] && !f[359] && f[384];
	assign leaf[3612] = f[325] && !f[357] && f[359] && !f[303];
	assign leaf[3613] = f[325] && !f[357] && f[359] && f[303];
	assign leaf[3614] = f[325] && f[357] && !f[268] && !f[214];
	assign leaf[3615] = f[325] && f[357] && !f[268] && f[214];
	assign leaf[3616] = f[325] && f[357] && f[268] && !f[490];
	assign leaf[3617] = f[325] && f[357] && f[268] && f[490];
	
	// Tree 237, Classifier 7, Iteration: 23
	assign leaf[3618] = !f[554] && !f[160] && !f[127] && !f[285];
	assign leaf[3619] = !f[554] && !f[160] && !f[127] && f[285];
	assign leaf[3620] = !f[554] && !f[160] && f[127] && !f[553];
	assign leaf[3621] = !f[554] && !f[160] && f[127] && f[553];
	assign leaf[3622] = !f[554] && f[160] && !f[152];
	assign leaf[3623] = !f[554] && f[160] && f[152];
	assign leaf[3624] = f[554] && !f[274] && !f[146] && !f[216];
	assign leaf[3625] = f[554] && !f[274] && !f[146] && f[216];
	assign leaf[3626] = f[554] && !f[274] && f[146];
	assign leaf[3627] = f[554] && f[274];
	
	// Tree 238, Classifier 8, Iteration: 23
	assign leaf[3628] = !f[301] && !f[330] && !f[271] && !f[300];
	assign leaf[3629] = !f[301] && !f[330] && !f[271] && f[300];
	assign leaf[3630] = !f[301] && !f[330] && f[271] && !f[242];
	assign leaf[3631] = !f[301] && !f[330] && f[271] && f[242];
	assign leaf[3632] = !f[301] && f[330] && !f[524] && !f[439];
	assign leaf[3633] = !f[301] && f[330] && !f[524] && f[439];
	assign leaf[3634] = !f[301] && f[330] && f[524];
	assign leaf[3635] = f[301] && !f[298] && !f[322] && !f[399];
	assign leaf[3636] = f[301] && !f[298] && !f[322] && f[399];
	assign leaf[3637] = f[301] && !f[298] && f[322] && !f[536];
	assign leaf[3638] = f[301] && !f[298] && f[322] && f[536];
	assign leaf[3639] = f[301] && f[298] && !f[458] && !f[459];
	assign leaf[3640] = f[301] && f[298] && !f[458] && f[459];
	assign leaf[3641] = f[301] && f[298] && f[458] && !f[243];
	assign leaf[3642] = f[301] && f[298] && f[458] && f[243];
	
	// Tree 239, Classifier 9, Iteration: 23
	assign leaf[3643] = !f[571] && !f[188] && !f[218] && !f[378];
	assign leaf[3644] = !f[571] && !f[188] && !f[218] && f[378];
	assign leaf[3645] = !f[571] && !f[188] && f[218] && !f[211];
	assign leaf[3646] = !f[571] && !f[188] && f[218] && f[211];
	assign leaf[3647] = !f[571] && f[188] && !f[383] && !f[545];
	assign leaf[3648] = !f[571] && f[188] && !f[383] && f[545];
	assign leaf[3649] = !f[571] && f[188] && f[383] && !f[574];
	assign leaf[3650] = !f[571] && f[188] && f[383] && f[574];
	assign leaf[3651] = f[571] && !f[213] && !f[425] && !f[574];
	assign leaf[3652] = f[571] && !f[213] && !f[425] && f[574];
	assign leaf[3653] = f[571] && !f[213] && f[425] && !f[240];
	assign leaf[3654] = f[571] && !f[213] && f[425] && f[240];
	assign leaf[3655] = f[571] && f[213] && !f[657] && !f[319];
	assign leaf[3656] = f[571] && f[213] && !f[657] && f[319];
	assign leaf[3657] = f[571] && f[213] && f[657] && !f[488];
	assign leaf[3658] = f[571] && f[213] && f[657] && f[488];
	
	// Tree 240, Classifier 0, Iteration: 24
	assign leaf[3659] = !f[663] && !f[406] && !f[688] && !f[398];
	assign leaf[3660] = !f[663] && !f[406] && !f[688] && f[398];
	assign leaf[3661] = !f[663] && !f[406] && f[688] && !f[656];
	assign leaf[3662] = !f[663] && !f[406] && f[688] && f[656];
	assign leaf[3663] = !f[663] && f[406] && !f[380] && !f[347];
	assign leaf[3664] = !f[663] && f[406] && !f[380] && f[347];
	assign leaf[3665] = !f[663] && f[406] && f[380] && !f[571];
	assign leaf[3666] = !f[663] && f[406] && f[380] && f[571];
	assign leaf[3667] = f[663] && !f[526] && !f[687] && !f[638];
	assign leaf[3668] = f[663] && !f[526] && !f[687] && f[638];
	assign leaf[3669] = f[663] && !f[526] && f[687] && !f[204];
	assign leaf[3670] = f[663] && !f[526] && f[687] && f[204];
	assign leaf[3671] = f[663] && f[526] && !f[347] && !f[402];
	assign leaf[3672] = f[663] && f[526] && !f[347] && f[402];
	assign leaf[3673] = f[663] && f[526] && f[347] && !f[572];
	assign leaf[3674] = f[663] && f[526] && f[347] && f[572];
	
	// Tree 241, Classifier 1, Iteration: 24
	assign leaf[3675] = !f[711] && !f[510] && !f[344] && !f[629];
	assign leaf[3676] = !f[711] && !f[510] && !f[344] && f[629];
	assign leaf[3677] = !f[711] && !f[510] && f[344] && !f[597];
	assign leaf[3678] = !f[711] && !f[510] && f[344] && f[597];
	assign leaf[3679] = !f[711] && f[510] && !f[484];
	assign leaf[3680] = !f[711] && f[510] && f[484] && !f[186];
	assign leaf[3681] = !f[711] && f[510] && f[484] && f[186];
	assign leaf[3682] = f[711] && !f[656];
	assign leaf[3683] = f[711] && f[656] && !f[710] && !f[294];
	assign leaf[3684] = f[711] && f[656] && !f[710] && f[294];
	assign leaf[3685] = f[711] && f[656] && f[710] && !f[354];
	assign leaf[3686] = f[711] && f[656] && f[710] && f[354];
	
	// Tree 242, Classifier 2, Iteration: 24
	assign leaf[3687] = !f[501] && !f[373] && !f[349] && !f[398];
	assign leaf[3688] = !f[501] && !f[373] && !f[349] && f[398];
	assign leaf[3689] = !f[501] && !f[373] && f[349] && !f[415];
	assign leaf[3690] = !f[501] && !f[373] && f[349] && f[415];
	assign leaf[3691] = !f[501] && f[373] && !f[426] && !f[547];
	assign leaf[3692] = !f[501] && f[373] && !f[426] && f[547];
	assign leaf[3693] = !f[501] && f[373] && f[426] && !f[290];
	assign leaf[3694] = !f[501] && f[373] && f[426] && f[290];
	assign leaf[3695] = f[501] && !f[370] && !f[654] && !f[264];
	assign leaf[3696] = f[501] && !f[370] && !f[654] && f[264];
	assign leaf[3697] = f[501] && !f[370] && f[654];
	assign leaf[3698] = f[501] && f[370];
	
	// Tree 243, Classifier 3, Iteration: 24
	assign leaf[3699] = !f[357] && !f[123] && !f[682] && !f[202];
	assign leaf[3700] = !f[357] && !f[123] && !f[682] && f[202];
	assign leaf[3701] = !f[357] && !f[123] && f[682] && !f[572];
	assign leaf[3702] = !f[357] && !f[123] && f[682] && f[572];
	assign leaf[3703] = !f[357] && f[123] && !f[234] && !f[260];
	assign leaf[3704] = !f[357] && f[123] && !f[234] && f[260];
	assign leaf[3705] = !f[357] && f[123] && f[234] && !f[147];
	assign leaf[3706] = !f[357] && f[123] && f[234] && f[147];
	assign leaf[3707] = f[357] && !f[355] && !f[488];
	assign leaf[3708] = f[357] && !f[355] && f[488] && !f[213];
	assign leaf[3709] = f[357] && !f[355] && f[488] && f[213];
	assign leaf[3710] = f[357] && f[355] && !f[399] && !f[239];
	assign leaf[3711] = f[357] && f[355] && !f[399] && f[239];
	assign leaf[3712] = f[357] && f[355] && f[399] && !f[160];
	assign leaf[3713] = f[357] && f[355] && f[399] && f[160];
	
	// Tree 244, Classifier 4, Iteration: 24
	assign leaf[3714] = !f[347] && !f[345] && !f[343] && !f[348];
	assign leaf[3715] = !f[347] && !f[345] && !f[343] && f[348];
	assign leaf[3716] = !f[347] && !f[345] && f[343] && !f[180];
	assign leaf[3717] = !f[347] && !f[345] && f[343] && f[180];
	assign leaf[3718] = !f[347] && f[345] && !f[454] && !f[236];
	assign leaf[3719] = !f[347] && f[345] && !f[454] && f[236];
	assign leaf[3720] = !f[347] && f[345] && f[454] && !f[320];
	assign leaf[3721] = !f[347] && f[345] && f[454] && f[320];
	assign leaf[3722] = f[347] && !f[408] && !f[324] && !f[382];
	assign leaf[3723] = f[347] && !f[408] && !f[324] && f[382];
	assign leaf[3724] = f[347] && !f[408] && f[324] && !f[407];
	assign leaf[3725] = f[347] && !f[408] && f[324] && f[407];
	assign leaf[3726] = f[347] && f[408] && !f[241] && !f[186];
	assign leaf[3727] = f[347] && f[408] && !f[241] && f[186];
	assign leaf[3728] = f[347] && f[408] && f[241] && !f[244];
	assign leaf[3729] = f[347] && f[408] && f[241] && f[244];
	
	// Tree 245, Classifier 5, Iteration: 24
	assign leaf[3730] = !f[380] && !f[325] && !f[411] && !f[242];
	assign leaf[3731] = !f[380] && !f[325] && !f[411] && f[242];
	assign leaf[3732] = !f[380] && !f[325] && f[411] && !f[520];
	assign leaf[3733] = !f[380] && !f[325] && f[411] && f[520];
	assign leaf[3734] = !f[380] && f[325] && !f[270] && !f[239];
	assign leaf[3735] = !f[380] && f[325] && !f[270] && f[239];
	assign leaf[3736] = !f[380] && f[325] && f[270] && !f[294];
	assign leaf[3737] = !f[380] && f[325] && f[270] && f[294];
	assign leaf[3738] = f[380] && !f[297] && !f[327] && !f[186];
	assign leaf[3739] = f[380] && !f[297] && !f[327] && f[186];
	assign leaf[3740] = f[380] && !f[297] && f[327] && !f[350];
	assign leaf[3741] = f[380] && !f[297] && f[327] && f[350];
	assign leaf[3742] = f[380] && f[297] && !f[274] && !f[295];
	assign leaf[3743] = f[380] && f[297] && !f[274] && f[295];
	assign leaf[3744] = f[380] && f[297] && f[274] && !f[354];
	assign leaf[3745] = f[380] && f[297] && f[274] && f[354];
	
	// Tree 246, Classifier 6, Iteration: 24
	assign leaf[3746] = !f[430] && !f[399] && !f[431] && !f[387];
	assign leaf[3747] = !f[430] && !f[399] && !f[431] && f[387];
	assign leaf[3748] = !f[430] && !f[399] && f[431] && !f[326];
	assign leaf[3749] = !f[430] && !f[399] && f[431] && f[326];
	assign leaf[3750] = !f[430] && f[399] && !f[434] && !f[432];
	assign leaf[3751] = !f[430] && f[399] && !f[434] && f[432];
	assign leaf[3752] = !f[430] && f[399] && f[434] && !f[546];
	assign leaf[3753] = !f[430] && f[399] && f[434] && f[546];
	assign leaf[3754] = f[430] && !f[486] && !f[432] && !f[300];
	assign leaf[3755] = f[430] && !f[486] && !f[432] && f[300];
	assign leaf[3756] = f[430] && !f[486] && f[432] && !f[487];
	assign leaf[3757] = f[430] && !f[486] && f[432] && f[487];
	assign leaf[3758] = f[430] && f[486] && !f[374] && !f[181];
	assign leaf[3759] = f[430] && f[486] && !f[374] && f[181];
	assign leaf[3760] = f[430] && f[486] && f[374] && !f[571];
	assign leaf[3761] = f[430] && f[486] && f[374] && f[571];
	
	// Tree 247, Classifier 7, Iteration: 24
	assign leaf[3762] = !f[298] && !f[347] && !f[687] && !f[685];
	assign leaf[3763] = !f[298] && !f[347] && !f[687] && f[685];
	assign leaf[3764] = !f[298] && !f[347] && f[687] && !f[574];
	assign leaf[3765] = !f[298] && !f[347] && f[687] && f[574];
	assign leaf[3766] = !f[298] && f[347] && !f[341] && !f[355];
	assign leaf[3767] = !f[298] && f[347] && !f[341] && f[355];
	assign leaf[3768] = !f[298] && f[347] && f[341] && !f[240];
	assign leaf[3769] = !f[298] && f[347] && f[341] && f[240];
	assign leaf[3770] = f[298] && !f[182] && !f[460] && !f[542];
	assign leaf[3771] = f[298] && !f[182] && !f[460] && f[542];
	assign leaf[3772] = f[298] && !f[182] && f[460] && !f[400];
	assign leaf[3773] = f[298] && !f[182] && f[460] && f[400];
	assign leaf[3774] = f[298] && f[182] && !f[633] && !f[576];
	assign leaf[3775] = f[298] && f[182] && !f[633] && f[576];
	assign leaf[3776] = f[298] && f[182] && f[633] && !f[716];
	assign leaf[3777] = f[298] && f[182] && f[633] && f[716];
	
	// Tree 248, Classifier 8, Iteration: 24
	assign leaf[3778] = !f[322] && !f[489] && !f[487] && !f[484];
	assign leaf[3779] = !f[322] && !f[489] && !f[487] && f[484];
	assign leaf[3780] = !f[322] && !f[489] && f[487] && !f[457];
	assign leaf[3781] = !f[322] && !f[489] && f[487] && f[457];
	assign leaf[3782] = !f[322] && f[489] && !f[376] && !f[402];
	assign leaf[3783] = !f[322] && f[489] && !f[376] && f[402];
	assign leaf[3784] = !f[322] && f[489] && f[376] && !f[430];
	assign leaf[3785] = !f[322] && f[489] && f[376] && f[430];
	assign leaf[3786] = f[322] && !f[239] && !f[155] && !f[602];
	assign leaf[3787] = f[322] && !f[239] && !f[155] && f[602];
	assign leaf[3788] = f[322] && !f[239] && f[155] && !f[293];
	assign leaf[3789] = f[322] && !f[239] && f[155] && f[293];
	assign leaf[3790] = f[322] && f[239] && !f[296] && !f[348];
	assign leaf[3791] = f[322] && f[239] && !f[296] && f[348];
	assign leaf[3792] = f[322] && f[239] && f[296] && !f[662];
	assign leaf[3793] = f[322] && f[239] && f[296] && f[662];
	
	// Tree 249, Classifier 9, Iteration: 24
	assign leaf[3794] = !f[571] && !f[443] && !f[569] && !f[176];
	assign leaf[3795] = !f[571] && !f[443] && !f[569] && f[176];
	assign leaf[3796] = !f[571] && !f[443] && f[569] && !f[486];
	assign leaf[3797] = !f[571] && !f[443] && f[569] && f[486];
	assign leaf[3798] = !f[571] && f[443] && !f[368] && !f[683];
	assign leaf[3799] = !f[571] && f[443] && !f[368] && f[683];
	assign leaf[3800] = !f[571] && f[443] && f[368];
	assign leaf[3801] = f[571] && !f[680] && !f[488] && !f[213];
	assign leaf[3802] = f[571] && !f[680] && !f[488] && f[213];
	assign leaf[3803] = f[571] && !f[680] && f[488] && !f[678];
	assign leaf[3804] = f[571] && !f[680] && f[488] && f[678];
	assign leaf[3805] = f[571] && f[680] && !f[207] && !f[215];
	assign leaf[3806] = f[571] && f[680] && !f[207] && f[215];
	assign leaf[3807] = f[571] && f[680] && f[207] && !f[345];
	assign leaf[3808] = f[571] && f[680] && f[207] && f[345];
	
	// Tree 250, Classifier 0, Iteration: 25
	assign leaf[3809] = !f[434] && !f[177] && !f[517] && !f[350];
	assign leaf[3810] = !f[434] && !f[177] && !f[517] && f[350];
	assign leaf[3811] = !f[434] && !f[177] && f[517] && !f[297];
	assign leaf[3812] = !f[434] && !f[177] && f[517] && f[297];
	assign leaf[3813] = !f[434] && f[177] && !f[397] && !f[596];
	assign leaf[3814] = !f[434] && f[177] && !f[397] && f[596];
	assign leaf[3815] = !f[434] && f[177] && f[397] && !f[633];
	assign leaf[3816] = !f[434] && f[177] && f[397] && f[633];
	assign leaf[3817] = f[434] && !f[569] && !f[161];
	assign leaf[3818] = f[434] && !f[569] && f[161];
	assign leaf[3819] = f[434] && f[569] && !f[428] && !f[601];
	assign leaf[3820] = f[434] && f[569] && !f[428] && f[601];
	assign leaf[3821] = f[434] && f[569] && f[428] && !f[431];
	assign leaf[3822] = f[434] && f[569] && f[428] && f[431];
	
	// Tree 251, Classifier 1, Iteration: 25
	assign leaf[3823] = !f[483] && !f[711] && !f[715] && !f[185];
	assign leaf[3824] = !f[483] && !f[711] && !f[715] && f[185];
	assign leaf[3825] = !f[483] && !f[711] && f[715] && !f[428];
	assign leaf[3826] = !f[483] && !f[711] && f[715] && f[428];
	assign leaf[3827] = !f[483] && f[711] && !f[265] && !f[460];
	assign leaf[3828] = !f[483] && f[711] && !f[265] && f[460];
	assign leaf[3829] = !f[483] && f[711] && f[265];
	assign leaf[3830] = f[483] && !f[651] && !f[656];
	assign leaf[3831] = f[483] && !f[651] && f[656] && !f[239];
	assign leaf[3832] = f[483] && !f[651] && f[656] && f[239];
	assign leaf[3833] = f[483] && f[651];
	
	// Tree 252, Classifier 2, Iteration: 25
	assign leaf[3834] = !f[352] && !f[566] && !f[407] && !f[371];
	assign leaf[3835] = !f[352] && !f[566] && !f[407] && f[371];
	assign leaf[3836] = !f[352] && !f[566] && f[407] && !f[512];
	assign leaf[3837] = !f[352] && !f[566] && f[407] && f[512];
	assign leaf[3838] = !f[352] && f[566] && !f[342] && !f[301];
	assign leaf[3839] = !f[352] && f[566] && !f[342] && f[301];
	assign leaf[3840] = !f[352] && f[566] && f[342] && !f[298];
	assign leaf[3841] = !f[352] && f[566] && f[342] && f[298];
	assign leaf[3842] = f[352] && !f[411] && !f[579] && !f[635];
	assign leaf[3843] = f[352] && !f[411] && !f[579] && f[635];
	assign leaf[3844] = f[352] && !f[411] && f[579] && !f[466];
	assign leaf[3845] = f[352] && !f[411] && f[579] && f[466];
	assign leaf[3846] = f[352] && f[411] && !f[388] && !f[445];
	assign leaf[3847] = f[352] && f[411] && !f[388] && f[445];
	assign leaf[3848] = f[352] && f[411] && f[388] && !f[234];
	assign leaf[3849] = f[352] && f[411] && f[388] && f[234];
	
	// Tree 253, Classifier 3, Iteration: 25
	assign leaf[3850] = !f[429] && !f[124] && !f[406] && !f[465];
	assign leaf[3851] = !f[429] && !f[124] && !f[406] && f[465];
	assign leaf[3852] = !f[429] && !f[124] && f[406] && !f[347];
	assign leaf[3853] = !f[429] && !f[124] && f[406] && f[347];
	assign leaf[3854] = !f[429] && f[124] && !f[207] && !f[233];
	assign leaf[3855] = !f[429] && f[124] && !f[207] && f[233];
	assign leaf[3856] = !f[429] && f[124] && f[207] && !f[210];
	assign leaf[3857] = !f[429] && f[124] && f[207] && f[210];
	assign leaf[3858] = f[429] && !f[511] && !f[404] && !f[554];
	assign leaf[3859] = f[429] && !f[511] && !f[404] && f[554];
	assign leaf[3860] = f[429] && !f[511] && f[404] && !f[344];
	assign leaf[3861] = f[429] && !f[511] && f[404] && f[344];
	assign leaf[3862] = f[429] && f[511] && !f[425] && !f[456];
	assign leaf[3863] = f[429] && f[511] && !f[425] && f[456];
	assign leaf[3864] = f[429] && f[511] && f[425] && !f[572];
	assign leaf[3865] = f[429] && f[511] && f[425] && f[572];
	
	// Tree 254, Classifier 4, Iteration: 25
	assign leaf[3866] = !f[346] && !f[207] && !f[263] && !f[571];
	assign leaf[3867] = !f[346] && !f[207] && !f[263] && f[571];
	assign leaf[3868] = !f[346] && !f[207] && f[263] && !f[260];
	assign leaf[3869] = !f[346] && !f[207] && f[263] && f[260];
	assign leaf[3870] = !f[346] && f[207] && !f[290] && !f[319];
	assign leaf[3871] = !f[346] && f[207] && !f[290] && f[319];
	assign leaf[3872] = !f[346] && f[207] && f[290] && !f[183];
	assign leaf[3873] = !f[346] && f[207] && f[290] && f[183];
	assign leaf[3874] = f[346] && !f[428] && !f[572] && !f[627];
	assign leaf[3875] = f[346] && !f[428] && !f[572] && f[627];
	assign leaf[3876] = f[346] && !f[428] && f[572] && !f[575];
	assign leaf[3877] = f[346] && !f[428] && f[572] && f[575];
	assign leaf[3878] = f[346] && f[428] && !f[214] && !f[211];
	assign leaf[3879] = f[346] && f[428] && !f[214] && f[211];
	assign leaf[3880] = f[346] && f[428] && f[214] && !f[273];
	assign leaf[3881] = f[346] && f[428] && f[214] && f[273];
	
	// Tree 255, Classifier 5, Iteration: 25
	assign leaf[3882] = !f[102] && !f[305] && !f[188] && !f[246];
	assign leaf[3883] = !f[102] && !f[305] && !f[188] && f[246];
	assign leaf[3884] = !f[102] && !f[305] && f[188] && !f[301];
	assign leaf[3885] = !f[102] && !f[305] && f[188] && f[301];
	assign leaf[3886] = !f[102] && f[305] && !f[384] && !f[183];
	assign leaf[3887] = !f[102] && f[305] && !f[384] && f[183];
	assign leaf[3888] = !f[102] && f[305] && f[384];
	assign leaf[3889] = f[102] && !f[207] && !f[324] && !f[571];
	assign leaf[3890] = f[102] && !f[207] && !f[324] && f[571];
	assign leaf[3891] = f[102] && !f[207] && f[324] && !f[348];
	assign leaf[3892] = f[102] && !f[207] && f[324] && f[348];
	assign leaf[3893] = f[102] && f[207] && !f[372] && !f[264];
	assign leaf[3894] = f[102] && f[207] && !f[372] && f[264];
	assign leaf[3895] = f[102] && f[207] && f[372];
	
	// Tree 256, Classifier 6, Iteration: 25
	assign leaf[3896] = !f[685] && !f[325] && !f[274] && !f[351];
	assign leaf[3897] = !f[685] && !f[325] && !f[274] && f[351];
	assign leaf[3898] = !f[685] && !f[325] && f[274] && !f[580];
	assign leaf[3899] = !f[685] && !f[325] && f[274] && f[580];
	assign leaf[3900] = !f[685] && f[325] && !f[357] && !f[359];
	assign leaf[3901] = !f[685] && f[325] && !f[357] && f[359];
	assign leaf[3902] = !f[685] && f[325] && f[357] && !f[410];
	assign leaf[3903] = !f[685] && f[325] && f[357] && f[410];
	assign leaf[3904] = f[685] && !f[599];
	assign leaf[3905] = f[685] && f[599] && !f[206] && !f[325];
	assign leaf[3906] = f[685] && f[599] && !f[206] && f[325];
	assign leaf[3907] = f[685] && f[599] && f[206];
	
	// Tree 257, Classifier 7, Iteration: 25
	assign leaf[3908] = !f[607] && !f[438] && !f[349] && !f[432];
	assign leaf[3909] = !f[607] && !f[438] && !f[349] && f[432];
	assign leaf[3910] = !f[607] && !f[438] && f[349] && !f[294];
	assign leaf[3911] = !f[607] && !f[438] && f[349] && f[294];
	assign leaf[3912] = !f[607] && f[438] && !f[540] && !f[372];
	assign leaf[3913] = !f[607] && f[438] && !f[540] && f[372];
	assign leaf[3914] = !f[607] && f[438] && f[540] && !f[233];
	assign leaf[3915] = !f[607] && f[438] && f[540] && f[233];
	assign leaf[3916] = f[607] && !f[435] && !f[180] && !f[319];
	assign leaf[3917] = f[607] && !f[435] && !f[180] && f[319];
	assign leaf[3918] = f[607] && !f[435] && f[180] && !f[173];
	assign leaf[3919] = f[607] && !f[435] && f[180] && f[173];
	assign leaf[3920] = f[607] && f[435] && !f[228] && !f[718];
	assign leaf[3921] = f[607] && f[435] && !f[228] && f[718];
	assign leaf[3922] = f[607] && f[435] && f[228] && !f[261];
	assign leaf[3923] = f[607] && f[435] && f[228] && f[261];
	
	// Tree 258, Classifier 8, Iteration: 25
	assign leaf[3924] = !f[287] && !f[468] && !f[357] && !f[410];
	assign leaf[3925] = !f[287] && !f[468] && !f[357] && f[410];
	assign leaf[3926] = !f[287] && !f[468] && f[357] && !f[327];
	assign leaf[3927] = !f[287] && !f[468] && f[357] && f[327];
	assign leaf[3928] = !f[287] && f[468] && !f[322] && !f[354];
	assign leaf[3929] = !f[287] && f[468] && !f[322] && f[354];
	assign leaf[3930] = !f[287] && f[468] && f[322] && !f[262];
	assign leaf[3931] = !f[287] && f[468] && f[322] && f[262];
	assign leaf[3932] = f[287] && !f[517] && !f[346] && !f[401];
	assign leaf[3933] = f[287] && !f[517] && !f[346] && f[401];
	assign leaf[3934] = f[287] && !f[517] && f[346] && !f[371];
	assign leaf[3935] = f[287] && !f[517] && f[346] && f[371];
	assign leaf[3936] = f[287] && f[517] && !f[514] && !f[682];
	assign leaf[3937] = f[287] && f[517] && !f[514] && f[682];
	assign leaf[3938] = f[287] && f[517] && f[514] && !f[343];
	assign leaf[3939] = f[287] && f[517] && f[514] && f[343];
	
	// Tree 259, Classifier 9, Iteration: 25
	assign leaf[3940] = !f[544] && !f[380] && !f[488] && !f[324];
	assign leaf[3941] = !f[544] && !f[380] && !f[488] && f[324];
	assign leaf[3942] = !f[544] && !f[380] && f[488] && !f[348];
	assign leaf[3943] = !f[544] && !f[380] && f[488] && f[348];
	assign leaf[3944] = !f[544] && f[380] && !f[467] && !f[412];
	assign leaf[3945] = !f[544] && f[380] && !f[467] && f[412];
	assign leaf[3946] = !f[544] && f[380] && f[467] && !f[356];
	assign leaf[3947] = !f[544] && f[380] && f[467] && f[356];
	assign leaf[3948] = f[544] && !f[629] && !f[488] && !f[273];
	assign leaf[3949] = f[544] && !f[629] && !f[488] && f[273];
	assign leaf[3950] = f[544] && !f[629] && f[488] && !f[399];
	assign leaf[3951] = f[544] && !f[629] && f[488] && f[399];
	assign leaf[3952] = f[544] && f[629] && !f[207] && !f[213];
	assign leaf[3953] = f[544] && f[629] && !f[207] && f[213];
	assign leaf[3954] = f[544] && f[629] && f[207] && !f[461];
	assign leaf[3955] = f[544] && f[629] && f[207] && f[461];
	
	// Tree 260, Classifier 0, Iteration: 26
	assign leaf[3956] = !f[542] && !f[510] && !f[512] && !f[471];
	assign leaf[3957] = !f[542] && !f[510] && !f[512] && f[471];
	assign leaf[3958] = !f[542] && !f[510] && f[512] && !f[654];
	assign leaf[3959] = !f[542] && !f[510] && f[512] && f[654];
	assign leaf[3960] = !f[542] && f[510] && !f[246] && !f[404];
	assign leaf[3961] = !f[542] && f[510] && !f[246] && f[404];
	assign leaf[3962] = !f[542] && f[510] && f[246] && !f[487];
	assign leaf[3963] = !f[542] && f[510] && f[246] && f[487];
	assign leaf[3964] = f[542] && !f[298] && !f[272] && !f[297];
	assign leaf[3965] = f[542] && !f[298] && !f[272] && f[297];
	assign leaf[3966] = f[542] && !f[298] && f[272] && !f[545];
	assign leaf[3967] = f[542] && !f[298] && f[272] && f[545];
	assign leaf[3968] = f[542] && f[298] && !f[430] && !f[415];
	assign leaf[3969] = f[542] && f[298] && !f[430] && f[415];
	assign leaf[3970] = f[542] && f[298] && f[430] && !f[383];
	assign leaf[3971] = f[542] && f[298] && f[430] && f[383];
	
	// Tree 261, Classifier 1, Iteration: 26
	assign leaf[3972] = !f[209] && !f[153] && !f[265] && !f[520];
	assign leaf[3973] = !f[209] && !f[153] && !f[265] && f[520];
	assign leaf[3974] = !f[209] && !f[153] && f[265] && !f[155];
	assign leaf[3975] = !f[209] && !f[153] && f[265] && f[155];
	assign leaf[3976] = !f[209] && f[153] && !f[488] && !f[99];
	assign leaf[3977] = !f[209] && f[153] && !f[488] && f[99];
	assign leaf[3978] = !f[209] && f[153] && f[488] && !f[539];
	assign leaf[3979] = !f[209] && f[153] && f[488] && f[539];
	assign leaf[3980] = f[209] && !f[266] && !f[378] && !f[128];
	assign leaf[3981] = f[209] && !f[266] && !f[378] && f[128];
	assign leaf[3982] = f[209] && !f[266] && f[378] && !f[268];
	assign leaf[3983] = f[209] && !f[266] && f[378] && f[268];
	assign leaf[3984] = f[209] && f[266] && !f[242] && !f[177];
	assign leaf[3985] = f[209] && f[266] && !f[242] && f[177];
	assign leaf[3986] = f[209] && f[266] && f[242] && !f[431];
	assign leaf[3987] = f[209] && f[266] && f[242] && f[431];
	
	// Tree 262, Classifier 2, Iteration: 26
	assign leaf[3988] = !f[152] && !f[497] && !f[580] && !f[415];
	assign leaf[3989] = !f[152] && !f[497] && !f[580] && f[415];
	assign leaf[3990] = !f[152] && !f[497] && f[580] && !f[260];
	assign leaf[3991] = !f[152] && !f[497] && f[580] && f[260];
	assign leaf[3992] = !f[152] && f[497] && !f[605] && !f[636];
	assign leaf[3993] = !f[152] && f[497] && !f[605] && f[636];
	assign leaf[3994] = !f[152] && f[497] && f[605] && !f[437];
	assign leaf[3995] = !f[152] && f[497] && f[605] && f[437];
	assign leaf[3996] = f[152] && !f[409] && !f[464] && !f[355];
	assign leaf[3997] = f[152] && !f[409] && !f[464] && f[355];
	assign leaf[3998] = f[152] && !f[409] && f[464] && !f[440];
	assign leaf[3999] = f[152] && !f[409] && f[464] && f[440];
	assign leaf[4000] = f[152] && f[409] && !f[519] && !f[438];
	assign leaf[4001] = f[152] && f[409] && !f[519] && f[438];
	assign leaf[4002] = f[152] && f[409] && f[519] && !f[609];
	assign leaf[4003] = f[152] && f[409] && f[519] && f[609];
	
	// Tree 263, Classifier 3, Iteration: 26
	assign leaf[4004] = !f[712] && !f[120] && !f[242] && !f[239];
	assign leaf[4005] = !f[712] && !f[120] && !f[242] && f[239];
	assign leaf[4006] = !f[712] && !f[120] && f[242] && !f[157];
	assign leaf[4007] = !f[712] && !f[120] && f[242] && f[157];
	assign leaf[4008] = !f[712] && f[120] && !f[632] && !f[293];
	assign leaf[4009] = !f[712] && f[120] && !f[632] && f[293];
	assign leaf[4010] = !f[712] && f[120] && f[632] && !f[235];
	assign leaf[4011] = !f[712] && f[120] && f[632] && f[235];
	assign leaf[4012] = f[712] && !f[601] && !f[376] && !f[435];
	assign leaf[4013] = f[712] && !f[601] && !f[376] && f[435];
	assign leaf[4014] = f[712] && !f[601] && f[376] && !f[232];
	assign leaf[4015] = f[712] && !f[601] && f[376] && f[232];
	assign leaf[4016] = f[712] && f[601] && !f[659] && !f[738];
	assign leaf[4017] = f[712] && f[601] && !f[659] && f[738];
	assign leaf[4018] = f[712] && f[601] && f[659] && !f[374];
	assign leaf[4019] = f[712] && f[601] && f[659] && f[374];
	
	// Tree 264, Classifier 4, Iteration: 26
	assign leaf[4020] = !f[740] && !f[409] && !f[438] && !f[577];
	assign leaf[4021] = !f[740] && !f[409] && !f[438] && f[577];
	assign leaf[4022] = !f[740] && !f[409] && f[438] && !f[248];
	assign leaf[4023] = !f[740] && !f[409] && f[438] && f[248];
	assign leaf[4024] = !f[740] && f[409] && !f[403] && !f[454];
	assign leaf[4025] = !f[740] && f[409] && !f[403] && f[454];
	assign leaf[4026] = !f[740] && f[409] && f[403] && !f[434];
	assign leaf[4027] = !f[740] && f[409] && f[403] && f[434];
	assign leaf[4028] = f[740] && !f[412];
	assign leaf[4029] = f[740] && f[412];
	
	// Tree 265, Classifier 5, Iteration: 26
	assign leaf[4030] = !f[485] && !f[541] && !f[379] && !f[409];
	assign leaf[4031] = !f[485] && !f[541] && !f[379] && f[409];
	assign leaf[4032] = !f[485] && !f[541] && f[379] && !f[324];
	assign leaf[4033] = !f[485] && !f[541] && f[379] && f[324];
	assign leaf[4034] = !f[485] && f[541] && !f[427] && !f[487];
	assign leaf[4035] = !f[485] && f[541] && !f[427] && f[487];
	assign leaf[4036] = !f[485] && f[541] && f[427] && !f[354];
	assign leaf[4037] = !f[485] && f[541] && f[427] && f[354];
	assign leaf[4038] = f[485] && !f[541] && !f[539] && !f[374];
	assign leaf[4039] = f[485] && !f[541] && !f[539] && f[374];
	assign leaf[4040] = f[485] && !f[541] && f[539] && !f[444];
	assign leaf[4041] = f[485] && !f[541] && f[539] && f[444];
	assign leaf[4042] = f[485] && f[541] && !f[430] && !f[428];
	assign leaf[4043] = f[485] && f[541] && !f[430] && f[428];
	assign leaf[4044] = f[485] && f[541] && f[430] && !f[276];
	assign leaf[4045] = f[485] && f[541] && f[430] && f[276];
	
	// Tree 266, Classifier 6, Iteration: 26
	assign leaf[4046] = !f[683] && !f[609] && !f[403] && !f[414];
	assign leaf[4047] = !f[683] && !f[609] && !f[403] && f[414];
	assign leaf[4048] = !f[683] && !f[609] && f[403] && !f[487];
	assign leaf[4049] = !f[683] && !f[609] && f[403] && f[487];
	assign leaf[4050] = !f[683] && f[609] && !f[455] && !f[487];
	assign leaf[4051] = !f[683] && f[609] && !f[455] && f[487];
	assign leaf[4052] = !f[683] && f[609] && f[455] && !f[638];
	assign leaf[4053] = !f[683] && f[609] && f[455] && f[638];
	assign leaf[4054] = f[683];
	
	// Tree 267, Classifier 7, Iteration: 26
	assign leaf[4055] = !f[159] && !f[124] && !f[582] && !f[349];
	assign leaf[4056] = !f[159] && !f[124] && !f[582] && f[349];
	assign leaf[4057] = !f[159] && !f[124] && f[582] && !f[722];
	assign leaf[4058] = !f[159] && !f[124] && f[582] && f[722];
	assign leaf[4059] = !f[159] && f[124] && !f[399];
	assign leaf[4060] = !f[159] && f[124] && f[399];
	assign leaf[4061] = f[159] && !f[205] && !f[679];
	assign leaf[4062] = f[159] && !f[205] && f[679] && !f[487];
	assign leaf[4063] = f[159] && !f[205] && f[679] && f[487];
	assign leaf[4064] = f[159] && f[205] && !f[297];
	assign leaf[4065] = f[159] && f[205] && f[297];
	
	// Tree 268, Classifier 8, Iteration: 26
	assign leaf[4066] = !f[469] && !f[287] && !f[274] && !f[330];
	assign leaf[4067] = !f[469] && !f[287] && !f[274] && f[330];
	assign leaf[4068] = !f[469] && !f[287] && f[274] && !f[677];
	assign leaf[4069] = !f[469] && !f[287] && f[274] && f[677];
	assign leaf[4070] = !f[469] && f[287] && !f[374] && !f[400];
	assign leaf[4071] = !f[469] && f[287] && !f[374] && f[400];
	assign leaf[4072] = !f[469] && f[287] && f[374] && !f[438];
	assign leaf[4073] = !f[469] && f[287] && f[374] && f[438];
	assign leaf[4074] = f[469] && !f[523] && !f[206] && !f[570];
	assign leaf[4075] = f[469] && !f[523] && !f[206] && f[570];
	assign leaf[4076] = f[469] && !f[523] && f[206] && !f[401];
	assign leaf[4077] = f[469] && !f[523] && f[206] && f[401];
	assign leaf[4078] = f[469] && f[523] && !f[569] && !f[161];
	assign leaf[4079] = f[469] && f[523] && !f[569] && f[161];
	assign leaf[4080] = f[469] && f[523] && f[569] && !f[414];
	assign leaf[4081] = f[469] && f[523] && f[569] && f[414];
	
	// Tree 269, Classifier 9, Iteration: 26
	assign leaf[4082] = !f[742] && !f[355] && !f[439] && !f[523];
	assign leaf[4083] = !f[742] && !f[355] && !f[439] && f[523];
	assign leaf[4084] = !f[742] && !f[355] && f[439] && !f[356];
	assign leaf[4085] = !f[742] && !f[355] && f[439] && f[356];
	assign leaf[4086] = !f[742] && f[355] && !f[213] && !f[318];
	assign leaf[4087] = !f[742] && f[355] && !f[213] && f[318];
	assign leaf[4088] = !f[742] && f[355] && f[213] && !f[566];
	assign leaf[4089] = !f[742] && f[355] && f[213] && f[566];
	assign leaf[4090] = f[742] && !f[323] && !f[488] && !f[406];
	assign leaf[4091] = f[742] && !f[323] && !f[488] && f[406];
	assign leaf[4092] = f[742] && !f[323] && f[488] && !f[546];
	assign leaf[4093] = f[742] && !f[323] && f[488] && f[546];
	assign leaf[4094] = f[742] && f[323] && !f[259] && !f[214];
	assign leaf[4095] = f[742] && f[323] && !f[259] && f[214];
	assign leaf[4096] = f[742] && f[323] && f[259] && !f[206];
	assign leaf[4097] = f[742] && f[323] && f[259] && f[206];
	
	// Tree 270, Classifier 0, Iteration: 27
	assign leaf[4098] = !f[378] && !f[571] && !f[654] && !f[415];
	assign leaf[4099] = !f[378] && !f[571] && !f[654] && f[415];
	assign leaf[4100] = !f[378] && !f[571] && f[654] && !f[455];
	assign leaf[4101] = !f[378] && !f[571] && f[654] && f[455];
	assign leaf[4102] = !f[378] && f[571] && !f[681] && !f[159];
	assign leaf[4103] = !f[378] && f[571] && !f[681] && f[159];
	assign leaf[4104] = !f[378] && f[571] && f[681] && !f[511];
	assign leaf[4105] = !f[378] && f[571] && f[681] && f[511];
	assign leaf[4106] = f[378] && !f[294] && !f[376] && !f[496];
	assign leaf[4107] = f[378] && !f[294] && !f[376] && f[496];
	assign leaf[4108] = f[378] && !f[294] && f[376] && !f[353];
	assign leaf[4109] = f[378] && !f[294] && f[376] && f[353];
	assign leaf[4110] = f[378] && f[294] && !f[245] && !f[438];
	assign leaf[4111] = f[378] && f[294] && !f[245] && f[438];
	assign leaf[4112] = f[378] && f[294] && f[245] && !f[352];
	assign leaf[4113] = f[378] && f[294] && f[245] && f[352];
	
	// Tree 271, Classifier 1, Iteration: 27
	assign leaf[4114] = !f[383] && !f[710] && !f[492] && !f[235];
	assign leaf[4115] = !f[383] && !f[710] && !f[492] && f[235];
	assign leaf[4116] = !f[383] && !f[710] && f[492] && !f[606];
	assign leaf[4117] = !f[383] && !f[710] && f[492] && f[606];
	assign leaf[4118] = !f[383] && f[710] && !f[238] && !f[601];
	assign leaf[4119] = !f[383] && f[710] && !f[238] && f[601];
	assign leaf[4120] = !f[383] && f[710] && f[238];
	assign leaf[4121] = f[383] && !f[218] && !f[681];
	assign leaf[4122] = f[383] && !f[218] && f[681];
	assign leaf[4123] = f[383] && f[218] && !f[325];
	assign leaf[4124] = f[383] && f[218] && f[325];
	
	// Tree 272, Classifier 2, Iteration: 27
	assign leaf[4125] = !f[372] && !f[347] && !f[397] && !f[679];
	assign leaf[4126] = !f[372] && !f[347] && !f[397] && f[679];
	assign leaf[4127] = !f[372] && !f[347] && f[397] && !f[313];
	assign leaf[4128] = !f[372] && !f[347] && f[397] && f[313];
	assign leaf[4129] = !f[372] && f[347] && !f[444] && !f[580];
	assign leaf[4130] = !f[372] && f[347] && !f[444] && f[580];
	assign leaf[4131] = !f[372] && f[347] && f[444] && !f[567];
	assign leaf[4132] = !f[372] && f[347] && f[444] && f[567];
	assign leaf[4133] = f[372] && !f[316] && !f[291] && !f[482];
	assign leaf[4134] = f[372] && !f[316] && !f[291] && f[482];
	assign leaf[4135] = f[372] && !f[316] && f[291] && !f[444];
	assign leaf[4136] = f[372] && !f[316] && f[291] && f[444];
	assign leaf[4137] = f[372] && f[316] && !f[400] && !f[515];
	assign leaf[4138] = f[372] && f[316] && !f[400] && f[515];
	assign leaf[4139] = f[372] && f[316] && f[400] && !f[652];
	assign leaf[4140] = f[372] && f[316] && f[400] && f[652];
	
	// Tree 273, Classifier 3, Iteration: 27
	assign leaf[4141] = !f[200] && !f[373] && !f[320] && !f[681];
	assign leaf[4142] = !f[200] && !f[373] && !f[320] && f[681];
	assign leaf[4143] = !f[200] && !f[373] && f[320] && !f[267];
	assign leaf[4144] = !f[200] && !f[373] && f[320] && f[267];
	assign leaf[4145] = !f[200] && f[373] && !f[321] && !f[345];
	assign leaf[4146] = !f[200] && f[373] && !f[321] && f[345];
	assign leaf[4147] = !f[200] && f[373] && f[321] && !f[256];
	assign leaf[4148] = !f[200] && f[373] && f[321] && f[256];
	assign leaf[4149] = f[200] && !f[314] && !f[298] && !f[410];
	assign leaf[4150] = f[200] && !f[314] && !f[298] && f[410];
	assign leaf[4151] = f[200] && !f[314] && f[298] && !f[547];
	assign leaf[4152] = f[200] && !f[314] && f[298] && f[547];
	assign leaf[4153] = f[200] && f[314];
	
	// Tree 274, Classifier 4, Iteration: 27
	assign leaf[4154] = !f[743] && !f[96] && !f[628] && !f[684];
	assign leaf[4155] = !f[743] && !f[96] && !f[628] && f[684];
	assign leaf[4156] = !f[743] && !f[96] && f[628] && !f[604];
	assign leaf[4157] = !f[743] && !f[96] && f[628] && f[604];
	assign leaf[4158] = !f[743] && f[96] && !f[574];
	assign leaf[4159] = !f[743] && f[96] && f[574];
	assign leaf[4160] = f[743] && !f[459] && !f[295];
	assign leaf[4161] = f[743] && !f[459] && f[295];
	assign leaf[4162] = f[743] && f[459];
	
	// Tree 275, Classifier 5, Iteration: 27
	assign leaf[4163] = !f[102] && !f[583] && !f[455] && !f[538];
	assign leaf[4164] = !f[102] && !f[583] && !f[455] && f[538];
	assign leaf[4165] = !f[102] && !f[583] && f[455] && !f[400];
	assign leaf[4166] = !f[102] && !f[583] && f[455] && f[400];
	assign leaf[4167] = !f[102] && f[583] && !f[399] && !f[406];
	assign leaf[4168] = !f[102] && f[583] && !f[399] && f[406];
	assign leaf[4169] = !f[102] && f[583] && f[399] && !f[482];
	assign leaf[4170] = !f[102] && f[583] && f[399] && f[482];
	assign leaf[4171] = f[102] && !f[352] && !f[159] && !f[211];
	assign leaf[4172] = f[102] && !f[352] && !f[159] && f[211];
	assign leaf[4173] = f[102] && !f[352] && f[159] && !f[381];
	assign leaf[4174] = f[102] && !f[352] && f[159] && f[381];
	assign leaf[4175] = f[102] && f[352] && !f[243] && !f[320];
	assign leaf[4176] = f[102] && f[352] && !f[243] && f[320];
	assign leaf[4177] = f[102] && f[352] && f[243];
	
	// Tree 276, Classifier 6, Iteration: 27
	assign leaf[4178] = !f[209] && !f[154] && !f[575] && !f[520];
	assign leaf[4179] = !f[209] && !f[154] && !f[575] && f[520];
	assign leaf[4180] = !f[209] && !f[154] && f[575] && !f[291];
	assign leaf[4181] = !f[209] && !f[154] && f[575] && f[291];
	assign leaf[4182] = !f[209] && f[154] && !f[416] && !f[183];
	assign leaf[4183] = !f[209] && f[154] && !f[416] && f[183];
	assign leaf[4184] = !f[209] && f[154] && f[416] && !f[383];
	assign leaf[4185] = !f[209] && f[154] && f[416] && f[383];
	assign leaf[4186] = f[209] && !f[128] && !f[99] && !f[130];
	assign leaf[4187] = f[209] && !f[128] && !f[99] && f[130];
	assign leaf[4188] = f[209] && !f[128] && f[99] && !f[410];
	assign leaf[4189] = f[209] && !f[128] && f[99] && f[410];
	assign leaf[4190] = f[209] && f[128] && !f[430] && !f[351];
	assign leaf[4191] = f[209] && f[128] && !f[430] && f[351];
	assign leaf[4192] = f[209] && f[128] && f[430] && !f[292];
	assign leaf[4193] = f[209] && f[128] && f[430] && f[292];
	
	// Tree 277, Classifier 7, Iteration: 27
	assign leaf[4194] = !f[581] && !f[566] && !f[128] && !f[240];
	assign leaf[4195] = !f[581] && !f[566] && !f[128] && f[240];
	assign leaf[4196] = !f[581] && !f[566] && f[128];
	assign leaf[4197] = !f[581] && f[566] && !f[620] && !f[178];
	assign leaf[4198] = !f[581] && f[566] && !f[620] && f[178];
	assign leaf[4199] = !f[581] && f[566] && f[620];
	assign leaf[4200] = f[581] && !f[292] && !f[127] && !f[721];
	assign leaf[4201] = f[581] && !f[292] && !f[127] && f[721];
	assign leaf[4202] = f[581] && !f[292] && f[127];
	assign leaf[4203] = f[581] && f[292] && !f[603] && !f[437];
	assign leaf[4204] = f[581] && f[292] && !f[603] && f[437];
	assign leaf[4205] = f[581] && f[292] && f[603] && !f[573];
	assign leaf[4206] = f[581] && f[292] && f[603] && f[573];
	
	// Tree 278, Classifier 8, Iteration: 27
	assign leaf[4207] = !f[441] && !f[314] && !f[437] && !f[406];
	assign leaf[4208] = !f[441] && !f[314] && !f[437] && f[406];
	assign leaf[4209] = !f[441] && !f[314] && f[437] && !f[152];
	assign leaf[4210] = !f[441] && !f[314] && f[437] && f[152];
	assign leaf[4211] = !f[441] && f[314] && !f[353] && !f[296];
	assign leaf[4212] = !f[441] && f[314] && !f[353] && f[296];
	assign leaf[4213] = !f[441] && f[314] && f[353] && !f[431];
	assign leaf[4214] = !f[441] && f[314] && f[353] && f[431];
	assign leaf[4215] = f[441] && !f[332] && !f[555] && !f[593];
	assign leaf[4216] = f[441] && !f[332] && !f[555] && f[593];
	assign leaf[4217] = f[441] && !f[332] && f[555] && !f[300];
	assign leaf[4218] = f[441] && !f[332] && f[555] && f[300];
	assign leaf[4219] = f[441] && f[332] && !f[549] && !f[187];
	assign leaf[4220] = f[441] && f[332] && !f[549] && f[187];
	assign leaf[4221] = f[441] && f[332] && f[549];
	
	// Tree 279, Classifier 9, Iteration: 27
	assign leaf[4222] = !f[201] && !f[694] && !f[517] && !f[543];
	assign leaf[4223] = !f[201] && !f[694] && !f[517] && f[543];
	assign leaf[4224] = !f[201] && !f[694] && f[517] && !f[658];
	assign leaf[4225] = !f[201] && !f[694] && f[517] && f[658];
	assign leaf[4226] = !f[201] && f[694] && !f[403] && !f[666];
	assign leaf[4227] = !f[201] && f[694] && !f[403] && f[666];
	assign leaf[4228] = !f[201] && f[694] && f[403] && !f[313];
	assign leaf[4229] = !f[201] && f[694] && f[403] && f[313];
	assign leaf[4230] = f[201] && !f[379] && !f[665];
	assign leaf[4231] = f[201] && !f[379] && f[665];
	assign leaf[4232] = f[201] && f[379];
	
	// Tree 280, Classifier 0, Iteration: 28
	assign leaf[4233] = !f[265] && !f[351] && !f[493] && !f[321];
	assign leaf[4234] = !f[265] && !f[351] && !f[493] && f[321];
	assign leaf[4235] = !f[265] && !f[351] && f[493] && !f[288];
	assign leaf[4236] = !f[265] && !f[351] && f[493] && f[288];
	assign leaf[4237] = !f[265] && f[351] && !f[216] && !f[347];
	assign leaf[4238] = !f[265] && f[351] && !f[216] && f[347];
	assign leaf[4239] = !f[265] && f[351] && f[216] && !f[353];
	assign leaf[4240] = !f[265] && f[351] && f[216] && f[353];
	assign leaf[4241] = f[265] && !f[416] && !f[347] && !f[469];
	assign leaf[4242] = f[265] && !f[416] && !f[347] && f[469];
	assign leaf[4243] = f[265] && !f[416] && f[347] && !f[635];
	assign leaf[4244] = f[265] && !f[416] && f[347] && f[635];
	assign leaf[4245] = f[265] && f[416] && !f[414];
	assign leaf[4246] = f[265] && f[416] && f[414] && !f[398];
	assign leaf[4247] = f[265] && f[416] && f[414] && f[398];
	
	// Tree 281, Classifier 1, Iteration: 28
	assign leaf[4248] = !f[485] && !f[274] && !f[710] && !f[686];
	assign leaf[4249] = !f[485] && !f[274] && !f[710] && f[686];
	assign leaf[4250] = !f[485] && !f[274] && f[710] && !f[210];
	assign leaf[4251] = !f[485] && !f[274] && f[710] && f[210];
	assign leaf[4252] = !f[485] && f[274];
	assign leaf[4253] = f[485] && !f[237] && !f[596] && !f[131];
	assign leaf[4254] = f[485] && !f[237] && !f[596] && f[131];
	assign leaf[4255] = f[485] && !f[237] && f[596] && !f[573];
	assign leaf[4256] = f[485] && !f[237] && f[596] && f[573];
	assign leaf[4257] = f[485] && f[237] && !f[347];
	assign leaf[4258] = f[485] && f[237] && f[347] && !f[607];
	assign leaf[4259] = f[485] && f[237] && f[347] && f[607];
	
	// Tree 282, Classifier 2, Iteration: 28
	assign leaf[4260] = !f[514] && !f[379] && !f[572] && !f[174];
	assign leaf[4261] = !f[514] && !f[379] && !f[572] && f[174];
	assign leaf[4262] = !f[514] && !f[379] && f[572] && !f[294];
	assign leaf[4263] = !f[514] && !f[379] && f[572] && f[294];
	assign leaf[4264] = !f[514] && f[379] && !f[517] && !f[427];
	assign leaf[4265] = !f[514] && f[379] && !f[517] && f[427];
	assign leaf[4266] = !f[514] && f[379] && f[517] && !f[215];
	assign leaf[4267] = !f[514] && f[379] && f[517] && f[215];
	assign leaf[4268] = f[514] && !f[460] && !f[624] && !f[404];
	assign leaf[4269] = f[514] && !f[460] && !f[624] && f[404];
	assign leaf[4270] = f[514] && !f[460] && f[624] && !f[545];
	assign leaf[4271] = f[514] && !f[460] && f[624] && f[545];
	assign leaf[4272] = f[514] && f[460] && !f[679] && !f[409];
	assign leaf[4273] = f[514] && f[460] && !f[679] && f[409];
	assign leaf[4274] = f[514] && f[460] && f[679] && !f[631];
	assign leaf[4275] = f[514] && f[460] && f[679] && f[631];
	
	// Tree 283, Classifier 3, Iteration: 28
	assign leaf[4276] = !f[429] && !f[98] && !f[467] && !f[571];
	assign leaf[4277] = !f[429] && !f[98] && !f[467] && f[571];
	assign leaf[4278] = !f[429] && !f[98] && f[467] && !f[407];
	assign leaf[4279] = !f[429] && !f[98] && f[467] && f[407];
	assign leaf[4280] = !f[429] && f[98] && !f[208] && !f[431];
	assign leaf[4281] = !f[429] && f[98] && !f[208] && f[431];
	assign leaf[4282] = !f[429] && f[98] && f[208] && !f[297];
	assign leaf[4283] = !f[429] && f[98] && f[208] && f[297];
	assign leaf[4284] = f[429] && !f[512] && !f[482] && !f[344];
	assign leaf[4285] = f[429] && !f[512] && !f[482] && f[344];
	assign leaf[4286] = f[429] && !f[512] && f[482] && !f[686];
	assign leaf[4287] = f[429] && !f[512] && f[482] && f[686];
	assign leaf[4288] = f[429] && f[512] && !f[453] && !f[201];
	assign leaf[4289] = f[429] && f[512] && !f[453] && f[201];
	assign leaf[4290] = f[429] && f[512] && f[453] && !f[432];
	assign leaf[4291] = f[429] && f[512] && f[453] && f[432];
	
	// Tree 284, Classifier 4, Iteration: 28
	assign leaf[4292] = !f[491] && !f[630] && !f[744] && !f[526];
	assign leaf[4293] = !f[491] && !f[630] && !f[744] && f[526];
	assign leaf[4294] = !f[491] && !f[630] && f[744];
	assign leaf[4295] = !f[491] && f[630] && !f[328] && !f[455];
	assign leaf[4296] = !f[491] && f[630] && !f[328] && f[455];
	assign leaf[4297] = !f[491] && f[630] && f[328] && !f[213];
	assign leaf[4298] = !f[491] && f[630] && f[328] && f[213];
	assign leaf[4299] = f[491] && !f[571] && !f[626] && !f[739];
	assign leaf[4300] = f[491] && !f[571] && !f[626] && f[739];
	assign leaf[4301] = f[491] && !f[571] && f[626] && !f[544];
	assign leaf[4302] = f[491] && !f[571] && f[626] && f[544];
	assign leaf[4303] = f[491] && f[571] && !f[186] && !f[654];
	assign leaf[4304] = f[491] && f[571] && !f[186] && f[654];
	assign leaf[4305] = f[491] && f[571] && f[186] && !f[497];
	assign leaf[4306] = f[491] && f[571] && f[186] && f[497];
	
	// Tree 285, Classifier 5, Iteration: 28
	assign leaf[4307] = !f[380] && !f[454] && !f[465] && !f[378];
	assign leaf[4308] = !f[380] && !f[454] && !f[465] && f[378];
	assign leaf[4309] = !f[380] && !f[454] && f[465] && !f[383];
	assign leaf[4310] = !f[380] && !f[454] && f[465] && f[383];
	assign leaf[4311] = !f[380] && f[454] && !f[407] && !f[399];
	assign leaf[4312] = !f[380] && f[454] && !f[407] && f[399];
	assign leaf[4313] = !f[380] && f[454] && f[407] && !f[440];
	assign leaf[4314] = !f[380] && f[454] && f[407] && f[440];
	assign leaf[4315] = f[380] && !f[434] && !f[297] && !f[294];
	assign leaf[4316] = f[380] && !f[434] && !f[297] && f[294];
	assign leaf[4317] = f[380] && !f[434] && f[297] && !f[154];
	assign leaf[4318] = f[380] && !f[434] && f[297] && f[154];
	assign leaf[4319] = f[380] && f[434] && !f[353] && !f[323];
	assign leaf[4320] = f[380] && f[434] && !f[353] && f[323];
	assign leaf[4321] = f[380] && f[434] && f[353] && !f[468];
	assign leaf[4322] = f[380] && f[434] && f[353] && f[468];
	
	// Tree 286, Classifier 6, Iteration: 28
	assign leaf[4323] = !f[686] && !f[623] && !f[163] && !f[269];
	assign leaf[4324] = !f[686] && !f[623] && !f[163] && f[269];
	assign leaf[4325] = !f[686] && !f[623] && f[163] && !f[597];
	assign leaf[4326] = !f[686] && !f[623] && f[163] && f[597];
	assign leaf[4327] = !f[686] && f[623] && !f[400] && !f[599];
	assign leaf[4328] = !f[686] && f[623] && !f[400] && f[599];
	assign leaf[4329] = !f[686] && f[623] && f[400] && !f[511];
	assign leaf[4330] = !f[686] && f[623] && f[400] && f[511];
	assign leaf[4331] = f[686] && !f[569];
	assign leaf[4332] = f[686] && f[569] && !f[234];
	assign leaf[4333] = f[686] && f[569] && f[234];
	
	// Tree 287, Classifier 7, Iteration: 28
	assign leaf[4334] = !f[124] && !f[161] && !f[527] && !f[266];
	assign leaf[4335] = !f[124] && !f[161] && !f[527] && f[266];
	assign leaf[4336] = !f[124] && !f[161] && f[527] && !f[511];
	assign leaf[4337] = !f[124] && !f[161] && f[527] && f[511];
	assign leaf[4338] = !f[124] && f[161] && !f[178];
	assign leaf[4339] = !f[124] && f[161] && f[178];
	assign leaf[4340] = f[124] && !f[427];
	assign leaf[4341] = f[124] && f[427];
	
	// Tree 288, Classifier 8, Iteration: 28
	assign leaf[4342] = !f[322] && !f[489] && !f[663] && !f[301];
	assign leaf[4343] = !f[322] && !f[489] && !f[663] && f[301];
	assign leaf[4344] = !f[322] && !f[489] && f[663] && !f[546];
	assign leaf[4345] = !f[322] && !f[489] && f[663] && f[546];
	assign leaf[4346] = !f[322] && f[489] && !f[485] && !f[659];
	assign leaf[4347] = !f[322] && f[489] && !f[485] && f[659];
	assign leaf[4348] = !f[322] && f[489] && f[485] && !f[493];
	assign leaf[4349] = !f[322] && f[489] && f[485] && f[493];
	assign leaf[4350] = f[322] && !f[546] && !f[264] && !f[290];
	assign leaf[4351] = f[322] && !f[546] && !f[264] && f[290];
	assign leaf[4352] = f[322] && !f[546] && f[264] && !f[238];
	assign leaf[4353] = f[322] && !f[546] && f[264] && f[238];
	assign leaf[4354] = f[322] && f[546] && !f[348] && !f[296];
	assign leaf[4355] = f[322] && f[546] && !f[348] && f[296];
	assign leaf[4356] = f[322] && f[546] && f[348] && !f[233];
	assign leaf[4357] = f[322] && f[546] && f[348] && f[233];
	
	// Tree 289, Classifier 9, Iteration: 28
	assign leaf[4358] = !f[594] && !f[129] && !f[149] && !f[379];
	assign leaf[4359] = !f[594] && !f[129] && !f[149] && f[379];
	assign leaf[4360] = !f[594] && !f[129] && f[149] && !f[258];
	assign leaf[4361] = !f[594] && !f[129] && f[149] && f[258];
	assign leaf[4362] = !f[594] && f[129] && !f[126];
	assign leaf[4363] = !f[594] && f[129] && f[126] && !f[292];
	assign leaf[4364] = !f[594] && f[129] && f[126] && f[292];
	assign leaf[4365] = f[594] && !f[551] && !f[181];
	assign leaf[4366] = f[594] && !f[551] && f[181] && !f[436];
	assign leaf[4367] = f[594] && !f[551] && f[181] && f[436];
	assign leaf[4368] = f[594] && f[551] && !f[399] && !f[211];
	assign leaf[4369] = f[594] && f[551] && !f[399] && f[211];
	assign leaf[4370] = f[594] && f[551] && f[399] && !f[466];
	assign leaf[4371] = f[594] && f[551] && f[399] && f[466];
	
	// Tree 290, Classifier 0, Iteration: 29
	assign leaf[4372] = !f[663] && !f[453] && !f[486] && !f[456];
	assign leaf[4373] = !f[663] && !f[453] && !f[486] && f[456];
	assign leaf[4374] = !f[663] && !f[453] && f[486] && !f[489];
	assign leaf[4375] = !f[663] && !f[453] && f[486] && f[489];
	assign leaf[4376] = !f[663] && f[453] && !f[303] && !f[329];
	assign leaf[4377] = !f[663] && f[453] && !f[303] && f[329];
	assign leaf[4378] = !f[663] && f[453] && f[303] && !f[150];
	assign leaf[4379] = !f[663] && f[453] && f[303] && f[150];
	assign leaf[4380] = f[663] && !f[498] && !f[630] && !f[689];
	assign leaf[4381] = f[663] && !f[498] && !f[630] && f[689];
	assign leaf[4382] = f[663] && !f[498] && f[630] && !f[604];
	assign leaf[4383] = f[663] && !f[498] && f[630] && f[604];
	assign leaf[4384] = f[663] && f[498] && !f[347] && !f[214];
	assign leaf[4385] = f[663] && f[498] && !f[347] && f[214];
	assign leaf[4386] = f[663] && f[498] && f[347] && !f[600];
	assign leaf[4387] = f[663] && f[498] && f[347] && f[600];
	
	// Tree 291, Classifier 1, Iteration: 29
	assign leaf[4388] = !f[440] && !f[301] && !f[520] && !f[207];
	assign leaf[4389] = !f[440] && !f[301] && !f[520] && f[207];
	assign leaf[4390] = !f[440] && !f[301] && f[520] && !f[606];
	assign leaf[4391] = !f[440] && !f[301] && f[520] && f[606];
	assign leaf[4392] = !f[440] && f[301] && !f[218];
	assign leaf[4393] = !f[440] && f[301] && f[218] && !f[239];
	assign leaf[4394] = !f[440] && f[301] && f[218] && f[239];
	assign leaf[4395] = f[440] && !f[300];
	assign leaf[4396] = f[440] && f[300];
	
	// Tree 292, Classifier 2, Iteration: 29
	assign leaf[4397] = !f[473] && !f[514] && !f[379] && !f[548];
	assign leaf[4398] = !f[473] && !f[514] && !f[379] && f[548];
	assign leaf[4399] = !f[473] && !f[514] && f[379] && !f[638];
	assign leaf[4400] = !f[473] && !f[514] && f[379] && f[638];
	assign leaf[4401] = !f[473] && f[514] && !f[433] && !f[353];
	assign leaf[4402] = !f[473] && f[514] && !f[433] && f[353];
	assign leaf[4403] = !f[473] && f[514] && f[433] && !f[651];
	assign leaf[4404] = !f[473] && f[514] && f[433] && f[651];
	assign leaf[4405] = f[473] && !f[343] && !f[354];
	assign leaf[4406] = f[473] && !f[343] && f[354];
	assign leaf[4407] = f[473] && f[343];
	
	// Tree 293, Classifier 3, Iteration: 29
	assign leaf[4408] = !f[678] && !f[147] && !f[318] && !f[292];
	assign leaf[4409] = !f[678] && !f[147] && !f[318] && f[292];
	assign leaf[4410] = !f[678] && !f[147] && f[318] && !f[293];
	assign leaf[4411] = !f[678] && !f[147] && f[318] && f[293];
	assign leaf[4412] = !f[678] && f[147] && !f[633] && !f[319];
	assign leaf[4413] = !f[678] && f[147] && !f[633] && f[319];
	assign leaf[4414] = !f[678] && f[147] && f[633] && !f[314];
	assign leaf[4415] = !f[678] && f[147] && f[633] && f[314];
	assign leaf[4416] = f[678] && !f[568] && !f[460] && !f[323];
	assign leaf[4417] = f[678] && !f[568] && !f[460] && f[323];
	assign leaf[4418] = f[678] && !f[568] && f[460] && !f[538];
	assign leaf[4419] = f[678] && !f[568] && f[460] && f[538];
	assign leaf[4420] = f[678] && f[568] && !f[514];
	assign leaf[4421] = f[678] && f[568] && f[514];
	
	// Tree 294, Classifier 4, Iteration: 29
	assign leaf[4422] = !f[286] && !f[594] && !f[348] && !f[345];
	assign leaf[4423] = !f[286] && !f[594] && !f[348] && f[345];
	assign leaf[4424] = !f[286] && !f[594] && f[348] && !f[381];
	assign leaf[4425] = !f[286] && !f[594] && f[348] && f[381];
	assign leaf[4426] = !f[286] && f[594] && !f[553] && !f[206];
	assign leaf[4427] = !f[286] && f[594] && !f[553] && f[206];
	assign leaf[4428] = !f[286] && f[594] && f[553];
	assign leaf[4429] = f[286] && !f[262] && !f[207] && !f[471];
	assign leaf[4430] = f[286] && !f[262] && !f[207] && f[471];
	assign leaf[4431] = f[286] && !f[262] && f[207] && !f[381];
	assign leaf[4432] = f[286] && !f[262] && f[207] && f[381];
	assign leaf[4433] = f[286] && f[262] && !f[218] && !f[396];
	assign leaf[4434] = f[286] && f[262] && !f[218] && f[396];
	assign leaf[4435] = f[286] && f[262] && f[218] && !f[412];
	assign leaf[4436] = f[286] && f[262] && f[218] && f[412];
	
	// Tree 295, Classifier 5, Iteration: 29
	assign leaf[4437] = !f[228] && !f[292] && !f[609] && !f[103];
	assign leaf[4438] = !f[228] && !f[292] && !f[609] && f[103];
	assign leaf[4439] = !f[228] && !f[292] && f[609] && !f[294];
	assign leaf[4440] = !f[228] && !f[292] && f[609] && f[294];
	assign leaf[4441] = !f[228] && f[292] && !f[235] && !f[125];
	assign leaf[4442] = !f[228] && f[292] && !f[235] && f[125];
	assign leaf[4443] = !f[228] && f[292] && f[235] && !f[457];
	assign leaf[4444] = !f[228] && f[292] && f[235] && f[457];
	assign leaf[4445] = f[228] && !f[172];
	assign leaf[4446] = f[228] && f[172];
	
	// Tree 296, Classifier 6, Iteration: 29
	assign leaf[4447] = !f[652] && !f[544] && !f[570] && !f[569];
	assign leaf[4448] = !f[652] && !f[544] && !f[570] && f[569];
	assign leaf[4449] = !f[652] && !f[544] && f[570] && !f[428];
	assign leaf[4450] = !f[652] && !f[544] && f[570] && f[428];
	assign leaf[4451] = !f[652] && f[544] && !f[236] && !f[153];
	assign leaf[4452] = !f[652] && f[544] && !f[236] && f[153];
	assign leaf[4453] = !f[652] && f[544] && f[236] && !f[322];
	assign leaf[4454] = !f[652] && f[544] && f[236] && f[322];
	assign leaf[4455] = f[652] && !f[133] && !f[498];
	assign leaf[4456] = f[652] && !f[133] && f[498];
	assign leaf[4457] = f[652] && f[133] && !f[292];
	assign leaf[4458] = f[652] && f[133] && f[292];
	
	// Tree 297, Classifier 7, Iteration: 29
	assign leaf[4459] = !f[744] && !f[577] && !f[662] && !f[207];
	assign leaf[4460] = !f[744] && !f[577] && !f[662] && f[207];
	assign leaf[4461] = !f[744] && !f[577] && f[662] && !f[178];
	assign leaf[4462] = !f[744] && !f[577] && f[662] && f[178];
	assign leaf[4463] = !f[744] && f[577] && !f[655] && !f[489];
	assign leaf[4464] = !f[744] && f[577] && !f[655] && f[489];
	assign leaf[4465] = !f[744] && f[577] && f[655] && !f[573];
	assign leaf[4466] = !f[744] && f[577] && f[655] && f[573];
	assign leaf[4467] = f[744] && !f[433] && !f[488] && !f[349];
	assign leaf[4468] = f[744] && !f[433] && !f[488] && f[349];
	assign leaf[4469] = f[744] && !f[433] && f[488] && !f[260];
	assign leaf[4470] = f[744] && !f[433] && f[488] && f[260];
	assign leaf[4471] = f[744] && f[433] && !f[440] && !f[294];
	assign leaf[4472] = f[744] && f[433] && !f[440] && f[294];
	assign leaf[4473] = f[744] && f[433] && f[440];
	
	// Tree 298, Classifier 8, Iteration: 29
	assign leaf[4474] = !f[261] && !f[374] && !f[292] && !f[266];
	assign leaf[4475] = !f[261] && !f[374] && !f[292] && f[266];
	assign leaf[4476] = !f[261] && !f[374] && f[292] && !f[238];
	assign leaf[4477] = !f[261] && !f[374] && f[292] && f[238];
	assign leaf[4478] = !f[261] && f[374] && !f[286] && !f[320];
	assign leaf[4479] = !f[261] && f[374] && !f[286] && f[320];
	assign leaf[4480] = !f[261] && f[374] && f[286] && !f[398];
	assign leaf[4481] = !f[261] && f[374] && f[286] && f[398];
	assign leaf[4482] = f[261] && !f[348] && !f[374] && !f[401];
	assign leaf[4483] = f[261] && !f[348] && !f[374] && f[401];
	assign leaf[4484] = f[261] && !f[348] && f[374] && !f[489];
	assign leaf[4485] = f[261] && !f[348] && f[374] && f[489];
	assign leaf[4486] = f[261] && f[348] && !f[372] && !f[235];
	assign leaf[4487] = f[261] && f[348] && !f[372] && f[235];
	assign leaf[4488] = f[261] && f[348] && f[372] && !f[434];
	assign leaf[4489] = f[261] && f[348] && f[372] && f[434];
	
	// Tree 299, Classifier 9, Iteration: 29
	assign leaf[4490] = !f[342] && !f[495] && !f[319] && !f[317];
	assign leaf[4491] = !f[342] && !f[495] && !f[319] && f[317];
	assign leaf[4492] = !f[342] && !f[495] && f[319] && !f[379];
	assign leaf[4493] = !f[342] && !f[495] && f[319] && f[379];
	assign leaf[4494] = !f[342] && f[495] && !f[664] && !f[344];
	assign leaf[4495] = !f[342] && f[495] && !f[664] && f[344];
	assign leaf[4496] = !f[342] && f[495] && f[664] && !f[607];
	assign leaf[4497] = !f[342] && f[495] && f[664] && f[607];
	assign leaf[4498] = f[342] && !f[345] && !f[385] && !f[213];
	assign leaf[4499] = f[342] && !f[345] && !f[385] && f[213];
	assign leaf[4500] = f[342] && !f[345] && f[385] && !f[343];
	assign leaf[4501] = f[342] && !f[345] && f[385] && f[343];
	assign leaf[4502] = f[342] && f[345] && !f[456] && !f[206];
	assign leaf[4503] = f[342] && f[345] && !f[456] && f[206];
	assign leaf[4504] = f[342] && f[345] && f[456] && !f[410];
	assign leaf[4505] = f[342] && f[345] && f[456] && f[410];
	
	// Tree 300, Classifier 0, Iteration: 30
	assign leaf[4506] = !f[444] && !f[213] && !f[240] && !f[326];
	assign leaf[4507] = !f[444] && !f[213] && !f[240] && f[326];
	assign leaf[4508] = !f[444] && !f[213] && f[240] && !f[542];
	assign leaf[4509] = !f[444] && !f[213] && f[240] && f[542];
	assign leaf[4510] = !f[444] && f[213] && !f[516] && !f[378];
	assign leaf[4511] = !f[444] && f[213] && !f[516] && f[378];
	assign leaf[4512] = !f[444] && f[213] && f[516] && !f[658];
	assign leaf[4513] = !f[444] && f[213] && f[516] && f[658];
	assign leaf[4514] = f[444] && !f[152] && !f[437] && !f[601];
	assign leaf[4515] = f[444] && !f[152] && !f[437] && f[601];
	assign leaf[4516] = f[444] && !f[152] && f[437];
	assign leaf[4517] = f[444] && f[152] && !f[302] && !f[299];
	assign leaf[4518] = f[444] && f[152] && !f[302] && f[299];
	assign leaf[4519] = f[444] && f[152] && f[302];
	
	// Tree 301, Classifier 1, Iteration: 30
	assign leaf[4520] = !f[439] && !f[272] && !f[294] && !f[182];
	assign leaf[4521] = !f[439] && !f[272] && !f[294] && f[182];
	assign leaf[4522] = !f[439] && !f[272] && f[294] && !f[189];
	assign leaf[4523] = !f[439] && !f[272] && f[294] && f[189];
	assign leaf[4524] = !f[439] && f[272] && !f[210] && !f[353];
	assign leaf[4525] = !f[439] && f[272] && !f[210] && f[353];
	assign leaf[4526] = !f[439] && f[272] && f[210] && !f[606];
	assign leaf[4527] = !f[439] && f[272] && f[210] && f[606];
	assign leaf[4528] = f[439] && !f[652];
	assign leaf[4529] = f[439] && f[652];
	
	// Tree 302, Classifier 2, Iteration: 30
	assign leaf[4530] = !f[682] && !f[713] && !f[372] && !f[351];
	assign leaf[4531] = !f[682] && !f[713] && !f[372] && f[351];
	assign leaf[4532] = !f[682] && !f[713] && f[372] && !f[316];
	assign leaf[4533] = !f[682] && !f[713] && f[372] && f[316];
	assign leaf[4534] = !f[682] && f[713] && !f[599];
	assign leaf[4535] = !f[682] && f[713] && f[599];
	assign leaf[4536] = f[682] && !f[180] && !f[605];
	assign leaf[4537] = f[682] && !f[180] && f[605];
	assign leaf[4538] = f[682] && f[180] && !f[431] && !f[406];
	assign leaf[4539] = f[682] && f[180] && !f[431] && f[406];
	assign leaf[4540] = f[682] && f[180] && f[431] && !f[541];
	assign leaf[4541] = f[682] && f[180] && f[431] && f[541];
	
	// Tree 303, Classifier 3, Iteration: 30
	assign leaf[4542] = !f[429] && !f[549] && !f[487] && !f[553];
	assign leaf[4543] = !f[429] && !f[549] && !f[487] && f[553];
	assign leaf[4544] = !f[429] && !f[549] && f[487] && !f[716];
	assign leaf[4545] = !f[429] && !f[549] && f[487] && f[716];
	assign leaf[4546] = !f[429] && f[549] && !f[712] && !f[263];
	assign leaf[4547] = !f[429] && f[549] && !f[712] && f[263];
	assign leaf[4548] = !f[429] && f[549] && f[712] && !f[320];
	assign leaf[4549] = !f[429] && f[549] && f[712] && f[320];
	assign leaf[4550] = f[429] && !f[433] && !f[516] && !f[482];
	assign leaf[4551] = f[429] && !f[433] && !f[516] && f[482];
	assign leaf[4552] = f[429] && !f[433] && f[516] && !f[464];
	assign leaf[4553] = f[429] && !f[433] && f[516] && f[464];
	assign leaf[4554] = f[429] && f[433] && !f[580] && !f[549];
	assign leaf[4555] = f[429] && f[433] && !f[580] && f[549];
	assign leaf[4556] = f[429] && f[433] && f[580] && !f[370];
	assign leaf[4557] = f[429] && f[433] && f[580] && f[370];
	
	// Tree 304, Classifier 4, Iteration: 30
	assign leaf[4558] = !f[745] && !f[399] && !f[375] && !f[373];
	assign leaf[4559] = !f[745] && !f[399] && !f[375] && f[373];
	assign leaf[4560] = !f[745] && !f[399] && f[375] && !f[601];
	assign leaf[4561] = !f[745] && !f[399] && f[375] && f[601];
	assign leaf[4562] = !f[745] && f[399] && !f[514] && !f[322];
	assign leaf[4563] = !f[745] && f[399] && !f[514] && f[322];
	assign leaf[4564] = !f[745] && f[399] && f[514] && !f[434];
	assign leaf[4565] = !f[745] && f[399] && f[514] && f[434];
	assign leaf[4566] = f[745] && !f[483];
	assign leaf[4567] = f[745] && f[483];
	
	// Tree 305, Classifier 5, Iteration: 30
	assign leaf[4568] = !f[684] && !f[600] && !f[603] && !f[440];
	assign leaf[4569] = !f[684] && !f[600] && !f[603] && f[440];
	assign leaf[4570] = !f[684] && !f[600] && f[603] && !f[628];
	assign leaf[4571] = !f[684] && !f[600] && f[603] && f[628];
	assign leaf[4572] = !f[684] && f[600] && !f[457] && !f[488];
	assign leaf[4573] = !f[684] && f[600] && !f[457] && f[488];
	assign leaf[4574] = !f[684] && f[600] && f[457] && !f[485];
	assign leaf[4575] = !f[684] && f[600] && f[457] && f[485];
	assign leaf[4576] = f[684] && !f[289] && !f[296] && !f[263];
	assign leaf[4577] = f[684] && !f[289] && !f[296] && f[263];
	assign leaf[4578] = f[684] && !f[289] && f[296] && !f[330];
	assign leaf[4579] = f[684] && !f[289] && f[296] && f[330];
	assign leaf[4580] = f[684] && f[289] && !f[578] && !f[373];
	assign leaf[4581] = f[684] && f[289] && !f[578] && f[373];
	assign leaf[4582] = f[684] && f[289] && f[578] && !f[401];
	assign leaf[4583] = f[684] && f[289] && f[578] && f[401];
	
	// Tree 306, Classifier 6, Iteration: 30
	assign leaf[4584] = !f[684] && !f[622] && !f[163] && !f[516];
	assign leaf[4585] = !f[684] && !f[622] && !f[163] && f[516];
	assign leaf[4586] = !f[684] && !f[622] && f[163] && !f[324];
	assign leaf[4587] = !f[684] && !f[622] && f[163] && f[324];
	assign leaf[4588] = !f[684] && f[622] && !f[498];
	assign leaf[4589] = !f[684] && f[622] && f[498];
	assign leaf[4590] = f[684] && !f[408] && !f[572];
	assign leaf[4591] = f[684] && !f[408] && f[572];
	assign leaf[4592] = f[684] && f[408];
	
	// Tree 307, Classifier 7, Iteration: 30
	assign leaf[4593] = !f[160] && !f[326] && !f[347] && !f[379];
	assign leaf[4594] = !f[160] && !f[326] && !f[347] && f[379];
	assign leaf[4595] = !f[160] && !f[326] && f[347] && !f[300];
	assign leaf[4596] = !f[160] && !f[326] && f[347] && f[300];
	assign leaf[4597] = !f[160] && f[326] && !f[433] && !f[488];
	assign leaf[4598] = !f[160] && f[326] && !f[433] && f[488];
	assign leaf[4599] = !f[160] && f[326] && f[433] && !f[489];
	assign leaf[4600] = !f[160] && f[326] && f[433] && f[489];
	assign leaf[4601] = f[160] && !f[687];
	assign leaf[4602] = f[160] && f[687];
	
	// Tree 308, Classifier 8, Iteration: 30
	assign leaf[4603] = !f[219] && !f[467] && !f[315] && !f[202];
	assign leaf[4604] = !f[219] && !f[467] && !f[315] && f[202];
	assign leaf[4605] = !f[219] && !f[467] && f[315] && !f[290];
	assign leaf[4606] = !f[219] && !f[467] && f[315] && f[290];
	assign leaf[4607] = !f[219] && f[467] && !f[521] && !f[638];
	assign leaf[4608] = !f[219] && f[467] && !f[521] && f[638];
	assign leaf[4609] = !f[219] && f[467] && f[521] && !f[637];
	assign leaf[4610] = !f[219] && f[467] && f[521] && f[637];
	assign leaf[4611] = f[219] && !f[458] && !f[655] && !f[685];
	assign leaf[4612] = f[219] && !f[458] && !f[655] && f[685];
	assign leaf[4613] = f[219] && !f[458] && f[655] && !f[346];
	assign leaf[4614] = f[219] && !f[458] && f[655] && f[346];
	assign leaf[4615] = f[219] && f[458] && !f[460] && !f[247];
	assign leaf[4616] = f[219] && f[458] && !f[460] && f[247];
	assign leaf[4617] = f[219] && f[458] && f[460] && !f[428];
	assign leaf[4618] = f[219] && f[458] && f[460] && f[428];
	
	// Tree 309, Classifier 9, Iteration: 30
	assign leaf[4619] = !f[161] && !f[572] && !f[188] && !f[209];
	assign leaf[4620] = !f[161] && !f[572] && !f[188] && f[209];
	assign leaf[4621] = !f[161] && !f[572] && f[188] && !f[601];
	assign leaf[4622] = !f[161] && !f[572] && f[188] && f[601];
	assign leaf[4623] = !f[161] && f[572] && !f[207] && !f[214];
	assign leaf[4624] = !f[161] && f[572] && !f[207] && f[214];
	assign leaf[4625] = !f[161] && f[572] && f[207] && !f[461];
	assign leaf[4626] = !f[161] && f[572] && f[207] && f[461];
	assign leaf[4627] = f[161] && !f[329];
	assign leaf[4628] = f[161] && f[329] && !f[601] && !f[319];
	assign leaf[4629] = f[161] && f[329] && !f[601] && f[319];
	assign leaf[4630] = f[161] && f[329] && f[601];
	
	// Tree 310, Classifier 0, Iteration: 31
	assign leaf[4631] = !f[204] && !f[664] && !f[415] && !f[241];
	assign leaf[4632] = !f[204] && !f[664] && !f[415] && f[241];
	assign leaf[4633] = !f[204] && !f[664] && f[415] && !f[436];
	assign leaf[4634] = !f[204] && !f[664] && f[415] && f[436];
	assign leaf[4635] = !f[204] && f[664] && !f[269];
	assign leaf[4636] = !f[204] && f[664] && f[269];
	assign leaf[4637] = f[204] && !f[398] && !f[399] && !f[272];
	assign leaf[4638] = f[204] && !f[398] && !f[399] && f[272];
	assign leaf[4639] = f[204] && !f[398] && f[399] && !f[513];
	assign leaf[4640] = f[204] && !f[398] && f[399] && f[513];
	assign leaf[4641] = f[204] && f[398] && !f[470] && !f[629];
	assign leaf[4642] = f[204] && f[398] && !f[470] && f[629];
	assign leaf[4643] = f[204] && f[398] && f[470] && !f[378];
	assign leaf[4644] = f[204] && f[398] && f[470] && f[378];
	
	// Tree 311, Classifier 1, Iteration: 31
	assign leaf[4645] = !f[456] && !f[490] && !f[629] && !f[658];
	assign leaf[4646] = !f[456] && !f[490] && !f[629] && f[658];
	assign leaf[4647] = !f[456] && !f[490] && f[629] && !f[378];
	assign leaf[4648] = !f[456] && !f[490] && f[629] && f[378];
	assign leaf[4649] = !f[456] && f[490] && !f[434] && !f[580];
	assign leaf[4650] = !f[456] && f[490] && !f[434] && f[580];
	assign leaf[4651] = !f[456] && f[490] && f[434] && !f[244];
	assign leaf[4652] = !f[456] && f[490] && f[434] && f[244];
	assign leaf[4653] = f[456] && !f[658] && !f[651];
	assign leaf[4654] = f[456] && !f[658] && f[651];
	assign leaf[4655] = f[456] && f[658] && !f[460];
	assign leaf[4656] = f[456] && f[658] && f[460];
	
	// Tree 312, Classifier 2, Iteration: 31
	assign leaf[4657] = !f[176] && !f[485] && !f[516] && !f[455];
	assign leaf[4658] = !f[176] && !f[485] && !f[516] && f[455];
	assign leaf[4659] = !f[176] && !f[485] && f[516] && !f[609];
	assign leaf[4660] = !f[176] && !f[485] && f[516] && f[609];
	assign leaf[4661] = !f[176] && f[485] && !f[432] && !f[595];
	assign leaf[4662] = !f[176] && f[485] && !f[432] && f[595];
	assign leaf[4663] = !f[176] && f[485] && f[432] && !f[685];
	assign leaf[4664] = !f[176] && f[485] && f[432] && f[685];
	assign leaf[4665] = f[176] && !f[551] && !f[691] && !f[341];
	assign leaf[4666] = f[176] && !f[551] && !f[691] && f[341];
	assign leaf[4667] = f[176] && !f[551] && f[691] && !f[610];
	assign leaf[4668] = f[176] && !f[551] && f[691] && f[610];
	assign leaf[4669] = f[176] && f[551] && !f[661] && !f[208];
	assign leaf[4670] = f[176] && f[551] && !f[661] && f[208];
	assign leaf[4671] = f[176] && f[551] && f[661] && !f[380];
	assign leaf[4672] = f[176] && f[551] && f[661] && f[380];
	
	// Tree 313, Classifier 3, Iteration: 31
	assign leaf[4673] = !f[399] && !f[536] && !f[551] && !f[125];
	assign leaf[4674] = !f[399] && !f[536] && !f[551] && f[125];
	assign leaf[4675] = !f[399] && !f[536] && f[551] && !f[238];
	assign leaf[4676] = !f[399] && !f[536] && f[551] && f[238];
	assign leaf[4677] = !f[399] && f[536] && !f[299] && !f[376];
	assign leaf[4678] = !f[399] && f[536] && !f[299] && f[376];
	assign leaf[4679] = !f[399] && f[536] && f[299] && !f[483];
	assign leaf[4680] = !f[399] && f[536] && f[299] && f[483];
	assign leaf[4681] = f[399] && !f[294] && !f[412] && !f[288];
	assign leaf[4682] = f[399] && !f[294] && !f[412] && f[288];
	assign leaf[4683] = f[399] && !f[294] && f[412] && !f[296];
	assign leaf[4684] = f[399] && !f[294] && f[412] && f[296];
	assign leaf[4685] = f[399] && f[294] && !f[288] && !f[526];
	assign leaf[4686] = f[399] && f[294] && !f[288] && f[526];
	assign leaf[4687] = f[399] && f[294] && f[288] && !f[516];
	assign leaf[4688] = f[399] && f[294] && f[288] && f[516];
	
	// Tree 314, Classifier 4, Iteration: 31
	assign leaf[4689] = !f[208] && !f[327] && !f[352] && !f[272];
	assign leaf[4690] = !f[208] && !f[327] && !f[352] && f[272];
	assign leaf[4691] = !f[208] && !f[327] && f[352] && !f[436];
	assign leaf[4692] = !f[208] && !f[327] && f[352] && f[436];
	assign leaf[4693] = !f[208] && f[327] && !f[241] && !f[296];
	assign leaf[4694] = !f[208] && f[327] && !f[241] && f[296];
	assign leaf[4695] = !f[208] && f[327] && f[241] && !f[467];
	assign leaf[4696] = !f[208] && f[327] && f[241] && f[467];
	assign leaf[4697] = f[208] && !f[184] && !f[239] && !f[243];
	assign leaf[4698] = f[208] && !f[184] && !f[239] && f[243];
	assign leaf[4699] = f[208] && !f[184] && f[239] && !f[234];
	assign leaf[4700] = f[208] && !f[184] && f[239] && f[234];
	assign leaf[4701] = f[208] && f[184] && !f[182] && !f[296];
	assign leaf[4702] = f[208] && f[184] && !f[182] && f[296];
	assign leaf[4703] = f[208] && f[184] && f[182] && !f[248];
	assign leaf[4704] = f[208] && f[184] && f[182] && f[248];
	
	// Tree 315, Classifier 5, Iteration: 31
	assign leaf[4705] = !f[277] && !f[628] && !f[548] && !f[332];
	assign leaf[4706] = !f[277] && !f[628] && !f[548] && f[332];
	assign leaf[4707] = !f[277] && !f[628] && f[548] && !f[683];
	assign leaf[4708] = !f[277] && !f[628] && f[548] && f[683];
	assign leaf[4709] = !f[277] && f[628] && !f[483] && !f[235];
	assign leaf[4710] = !f[277] && f[628] && !f[483] && f[235];
	assign leaf[4711] = !f[277] && f[628] && f[483] && !f[400];
	assign leaf[4712] = !f[277] && f[628] && f[483] && f[400];
	assign leaf[4713] = f[277] && !f[274];
	assign leaf[4714] = f[277] && f[274] && !f[651];
	assign leaf[4715] = f[277] && f[274] && f[651];
	
	// Tree 316, Classifier 6, Iteration: 31
	assign leaf[4716] = !f[602] && !f[547] && !f[630] && !f[164];
	assign leaf[4717] = !f[602] && !f[547] && !f[630] && f[164];
	assign leaf[4718] = !f[602] && !f[547] && f[630] && !f[206];
	assign leaf[4719] = !f[602] && !f[547] && f[630] && f[206];
	assign leaf[4720] = !f[602] && f[547] && !f[236] && !f[155];
	assign leaf[4721] = !f[602] && f[547] && !f[236] && f[155];
	assign leaf[4722] = !f[602] && f[547] && f[236] && !f[383];
	assign leaf[4723] = !f[602] && f[547] && f[236] && f[383];
	assign leaf[4724] = f[602] && !f[400] && !f[459] && !f[359];
	assign leaf[4725] = f[602] && !f[400] && !f[459] && f[359];
	assign leaf[4726] = f[602] && !f[400] && f[459] && !f[326];
	assign leaf[4727] = f[602] && !f[400] && f[459] && f[326];
	assign leaf[4728] = f[602] && f[400] && !f[382] && !f[483];
	assign leaf[4729] = f[602] && f[400] && !f[382] && f[483];
	assign leaf[4730] = f[602] && f[400] && f[382] && !f[441];
	assign leaf[4731] = f[602] && f[400] && f[382] && f[441];
	
	// Tree 317, Classifier 7, Iteration: 31
	assign leaf[4732] = !f[677] && !f[595] && !f[542] && !f[294];
	assign leaf[4733] = !f[677] && !f[595] && !f[542] && f[294];
	assign leaf[4734] = !f[677] && !f[595] && f[542] && !f[241];
	assign leaf[4735] = !f[677] && !f[595] && f[542] && f[241];
	assign leaf[4736] = !f[677] && f[595] && !f[292] && !f[681];
	assign leaf[4737] = !f[677] && f[595] && !f[292] && f[681];
	assign leaf[4738] = !f[677] && f[595] && f[292];
	assign leaf[4739] = f[677] && !f[682] && !f[516];
	assign leaf[4740] = f[677] && !f[682] && f[516] && !f[234];
	assign leaf[4741] = f[677] && !f[682] && f[516] && f[234];
	assign leaf[4742] = f[677] && f[682];
	
	// Tree 318, Classifier 8, Iteration: 31
	assign leaf[4743] = !f[439] && !f[525] && !f[542] && !f[512];
	assign leaf[4744] = !f[439] && !f[525] && !f[542] && f[512];
	assign leaf[4745] = !f[439] && !f[525] && f[542] && !f[544];
	assign leaf[4746] = !f[439] && !f[525] && f[542] && f[544];
	assign leaf[4747] = !f[439] && f[525] && !f[637] && !f[383];
	assign leaf[4748] = !f[439] && f[525] && !f[637] && f[383];
	assign leaf[4749] = !f[439] && f[525] && f[637] && !f[377];
	assign leaf[4750] = !f[439] && f[525] && f[637] && f[377];
	assign leaf[4751] = f[439] && !f[521] && !f[271] && !f[217];
	assign leaf[4752] = f[439] && !f[521] && !f[271] && f[217];
	assign leaf[4753] = f[439] && !f[521] && f[271] && !f[298];
	assign leaf[4754] = f[439] && !f[521] && f[271] && f[298];
	assign leaf[4755] = f[439] && f[521] && !f[594] && !f[153];
	assign leaf[4756] = f[439] && f[521] && !f[594] && f[153];
	assign leaf[4757] = f[439] && f[521] && f[594] && !f[457];
	assign leaf[4758] = f[439] && f[521] && f[594] && f[457];
	
	// Tree 319, Classifier 9, Iteration: 31
	assign leaf[4759] = !f[631] && !f[715] && !f[566] && !f[350];
	assign leaf[4760] = !f[631] && !f[715] && !f[566] && f[350];
	assign leaf[4761] = !f[631] && !f[715] && f[566] && !f[606];
	assign leaf[4762] = !f[631] && !f[715] && f[566] && f[606];
	assign leaf[4763] = !f[631] && f[715] && !f[381] && !f[294];
	assign leaf[4764] = !f[631] && f[715] && !f[381] && f[294];
	assign leaf[4765] = !f[631] && f[715] && f[381] && !f[743];
	assign leaf[4766] = !f[631] && f[715] && f[381] && f[743];
	assign leaf[4767] = f[631] && !f[545] && !f[209] && !f[742];
	assign leaf[4768] = f[631] && !f[545] && !f[209] && f[742];
	assign leaf[4769] = f[631] && !f[545] && f[209] && !f[237];
	assign leaf[4770] = f[631] && !f[545] && f[209] && f[237];
	assign leaf[4771] = f[631] && f[545] && !f[485] && !f[489];
	assign leaf[4772] = f[631] && f[545] && !f[485] && f[489];
	assign leaf[4773] = f[631] && f[545] && f[485] && !f[576];
	assign leaf[4774] = f[631] && f[545] && f[485] && f[576];
	
	// Tree 320, Classifier 0, Iteration: 32
	assign leaf[4775] = !f[688] && !f[103] && !f[663] && !f[406];
	assign leaf[4776] = !f[688] && !f[103] && !f[663] && f[406];
	assign leaf[4777] = !f[688] && !f[103] && f[663] && !f[659];
	assign leaf[4778] = !f[688] && !f[103] && f[663] && f[659];
	assign leaf[4779] = !f[688] && f[103] && !f[517] && !f[301];
	assign leaf[4780] = !f[688] && f[103] && !f[517] && f[301];
	assign leaf[4781] = !f[688] && f[103] && f[517] && !f[604];
	assign leaf[4782] = !f[688] && f[103] && f[517] && f[604];
	assign leaf[4783] = f[688] && !f[657] && !f[574] && !f[156];
	assign leaf[4784] = f[688] && !f[657] && !f[574] && f[156];
	assign leaf[4785] = f[688] && !f[657] && f[574];
	assign leaf[4786] = f[688] && f[657] && !f[571] && !f[347];
	assign leaf[4787] = f[688] && f[657] && !f[571] && f[347];
	assign leaf[4788] = f[688] && f[657] && f[571] && !f[523];
	assign leaf[4789] = f[688] && f[657] && f[571] && f[523];
	
	// Tree 321, Classifier 1, Iteration: 32
	assign leaf[4790] = !f[316] && !f[711] && !f[540] && !f[515];
	assign leaf[4791] = !f[316] && !f[711] && !f[540] && f[515];
	assign leaf[4792] = !f[316] && !f[711] && f[540] && !f[542];
	assign leaf[4793] = !f[316] && !f[711] && f[540] && f[542];
	assign leaf[4794] = !f[316] && f[711];
	assign leaf[4795] = f[316] && !f[127] && !f[159] && !f[151];
	assign leaf[4796] = f[316] && !f[127] && !f[159] && f[151];
	assign leaf[4797] = f[316] && !f[127] && f[159];
	assign leaf[4798] = f[316] && f[127] && !f[265];
	assign leaf[4799] = f[316] && f[127] && f[265];
	
	// Tree 322, Classifier 2, Iteration: 32
	assign leaf[4800] = !f[121] && !f[545] && !f[509] && !f[417];
	assign leaf[4801] = !f[121] && !f[545] && !f[509] && f[417];
	assign leaf[4802] = !f[121] && !f[545] && f[509] && !f[434];
	assign leaf[4803] = !f[121] && !f[545] && f[509] && f[434];
	assign leaf[4804] = !f[121] && f[545] && !f[634] && !f[551];
	assign leaf[4805] = !f[121] && f[545] && !f[634] && f[551];
	assign leaf[4806] = !f[121] && f[545] && f[634] && !f[495];
	assign leaf[4807] = !f[121] && f[545] && f[634] && f[495];
	assign leaf[4808] = f[121] && !f[232] && !f[290] && !f[605];
	assign leaf[4809] = f[121] && !f[232] && !f[290] && f[605];
	assign leaf[4810] = f[121] && !f[232] && f[290];
	assign leaf[4811] = f[121] && f[232] && !f[496] && !f[181];
	assign leaf[4812] = f[121] && f[232] && !f[496] && f[181];
	assign leaf[4813] = f[121] && f[232] && f[496] && !f[633];
	assign leaf[4814] = f[121] && f[232] && f[496] && f[633];
	
	// Tree 323, Classifier 3, Iteration: 32
	assign leaf[4815] = !f[370] && !f[346] && !f[320] && !f[372];
	assign leaf[4816] = !f[370] && !f[346] && !f[320] && f[372];
	assign leaf[4817] = !f[370] && !f[346] && f[320] && !f[292];
	assign leaf[4818] = !f[370] && !f[346] && f[320] && f[292];
	assign leaf[4819] = !f[370] && f[346] && !f[321] && !f[375];
	assign leaf[4820] = !f[370] && f[346] && !f[321] && f[375];
	assign leaf[4821] = !f[370] && f[346] && f[321] && !f[263];
	assign leaf[4822] = !f[370] && f[346] && f[321] && f[263];
	assign leaf[4823] = f[370] && !f[711] && !f[314] && !f[377];
	assign leaf[4824] = f[370] && !f[711] && !f[314] && f[377];
	assign leaf[4825] = f[370] && !f[711] && f[314] && !f[284];
	assign leaf[4826] = f[370] && !f[711] && f[314] && f[284];
	assign leaf[4827] = f[370] && f[711];
	
	// Tree 324, Classifier 4, Iteration: 32
	assign leaf[4828] = !f[219] && !f[286] && !f[600] && !f[655];
	assign leaf[4829] = !f[219] && !f[286] && !f[600] && f[655];
	assign leaf[4830] = !f[219] && !f[286] && f[600] && !f[576];
	assign leaf[4831] = !f[219] && !f[286] && f[600] && f[576];
	assign leaf[4832] = !f[219] && f[286] && !f[234] && !f[290];
	assign leaf[4833] = !f[219] && f[286] && !f[234] && f[290];
	assign leaf[4834] = !f[219] && f[286] && f[234] && !f[329];
	assign leaf[4835] = !f[219] && f[286] && f[234] && f[329];
	assign leaf[4836] = f[219] && !f[242] && !f[323] && !f[187];
	assign leaf[4837] = f[219] && !f[242] && !f[323] && f[187];
	assign leaf[4838] = f[219] && !f[242] && f[323] && !f[487];
	assign leaf[4839] = f[219] && !f[242] && f[323] && f[487];
	assign leaf[4840] = f[219] && f[242] && !f[240] && !f[655];
	assign leaf[4841] = f[219] && f[242] && !f[240] && f[655];
	assign leaf[4842] = f[219] && f[242] && f[240];
	
	// Tree 325, Classifier 5, Iteration: 32
	assign leaf[4843] = !f[490] && !f[103] && !f[609] && !f[263];
	assign leaf[4844] = !f[490] && !f[103] && !f[609] && f[263];
	assign leaf[4845] = !f[490] && !f[103] && f[609] && !f[287];
	assign leaf[4846] = !f[490] && !f[103] && f[609] && f[287];
	assign leaf[4847] = !f[490] && f[103] && !f[405] && !f[577];
	assign leaf[4848] = !f[490] && f[103] && !f[405] && f[577];
	assign leaf[4849] = !f[490] && f[103] && f[405] && !f[573];
	assign leaf[4850] = !f[490] && f[103] && f[405] && f[573];
	assign leaf[4851] = f[490] && !f[304] && !f[354] && !f[324];
	assign leaf[4852] = f[490] && !f[304] && !f[354] && f[324];
	assign leaf[4853] = f[490] && !f[304] && f[354] && !f[323];
	assign leaf[4854] = f[490] && !f[304] && f[354] && f[323];
	assign leaf[4855] = f[490] && f[304] && !f[300];
	assign leaf[4856] = f[490] && f[304] && f[300] && !f[599];
	assign leaf[4857] = f[490] && f[304] && f[300] && f[599];
	
	// Tree 326, Classifier 6, Iteration: 32
	assign leaf[4858] = !f[522] && !f[409] && !f[519] && !f[525];
	assign leaf[4859] = !f[522] && !f[409] && !f[519] && f[525];
	assign leaf[4860] = !f[522] && !f[409] && f[519] && !f[209];
	assign leaf[4861] = !f[522] && !f[409] && f[519] && f[209];
	assign leaf[4862] = !f[522] && f[409] && !f[525] && !f[319];
	assign leaf[4863] = !f[522] && f[409] && !f[525] && f[319];
	assign leaf[4864] = !f[522] && f[409] && f[525] && !f[322];
	assign leaf[4865] = !f[522] && f[409] && f[525] && f[322];
	assign leaf[4866] = f[522] && !f[402] && !f[387] && !f[212];
	assign leaf[4867] = f[522] && !f[402] && !f[387] && f[212];
	assign leaf[4868] = f[522] && !f[402] && f[387] && !f[264];
	assign leaf[4869] = f[522] && !f[402] && f[387] && f[264];
	assign leaf[4870] = f[522] && f[402] && !f[178] && !f[301];
	assign leaf[4871] = f[522] && f[402] && !f[178] && f[301];
	assign leaf[4872] = f[522] && f[402] && f[178] && !f[210];
	assign leaf[4873] = f[522] && f[402] && f[178] && f[210];
	
	// Tree 327, Classifier 7, Iteration: 32
	assign leaf[4874] = !f[609] && !f[549] && !f[206] && !f[260];
	assign leaf[4875] = !f[609] && !f[549] && !f[206] && f[260];
	assign leaf[4876] = !f[609] && !f[549] && f[206] && !f[634];
	assign leaf[4877] = !f[609] && !f[549] && f[206] && f[634];
	assign leaf[4878] = !f[609] && f[549] && !f[434] && !f[626];
	assign leaf[4879] = !f[609] && f[549] && !f[434] && f[626];
	assign leaf[4880] = !f[609] && f[549] && f[434] && !f[202];
	assign leaf[4881] = !f[609] && f[549] && f[434] && f[202];
	assign leaf[4882] = f[609] && !f[319] && !f[720];
	assign leaf[4883] = f[609] && !f[319] && f[720] && !f[294];
	assign leaf[4884] = f[609] && !f[319] && f[720] && f[294];
	assign leaf[4885] = f[609] && f[319] && !f[262];
	assign leaf[4886] = f[609] && f[319] && f[262] && !f[397];
	assign leaf[4887] = f[609] && f[319] && f[262] && f[397];
	
	// Tree 328, Classifier 8, Iteration: 32
	assign leaf[4888] = !f[441] && !f[341] && !f[357] && !f[410];
	assign leaf[4889] = !f[441] && !f[341] && !f[357] && f[410];
	assign leaf[4890] = !f[441] && !f[341] && f[357] && !f[328];
	assign leaf[4891] = !f[441] && !f[341] && f[357] && f[328];
	assign leaf[4892] = !f[441] && f[341] && !f[315] && !f[430];
	assign leaf[4893] = !f[441] && f[341] && !f[315] && f[430];
	assign leaf[4894] = !f[441] && f[341] && f[315] && !f[435];
	assign leaf[4895] = !f[441] && f[341] && f[315] && f[435];
	assign leaf[4896] = f[441] && !f[595] && !f[523] && !f[633];
	assign leaf[4897] = f[441] && !f[595] && !f[523] && f[633];
	assign leaf[4898] = f[441] && !f[595] && f[523] && !f[691];
	assign leaf[4899] = f[441] && !f[595] && f[523] && f[691];
	assign leaf[4900] = f[441] && f[595] && !f[496] && !f[510];
	assign leaf[4901] = f[441] && f[595] && !f[496] && f[510];
	assign leaf[4902] = f[441] && f[595] && f[496] && !f[456];
	assign leaf[4903] = f[441] && f[595] && f[496] && f[456];
	
	// Tree 329, Classifier 9, Iteration: 32
	assign leaf[4904] = !f[693] && !f[608] && !f[351] && !f[385];
	assign leaf[4905] = !f[693] && !f[608] && !f[351] && f[385];
	assign leaf[4906] = !f[693] && !f[608] && f[351] && !f[461];
	assign leaf[4907] = !f[693] && !f[608] && f[351] && f[461];
	assign leaf[4908] = !f[693] && f[608] && !f[692] && !f[330];
	assign leaf[4909] = !f[693] && f[608] && !f[692] && f[330];
	assign leaf[4910] = !f[693] && f[608] && f[692] && !f[318];
	assign leaf[4911] = !f[693] && f[608] && f[692] && f[318];
	assign leaf[4912] = f[693] && !f[229] && !f[320] && !f[203];
	assign leaf[4913] = f[693] && !f[229] && !f[320] && f[203];
	assign leaf[4914] = f[693] && !f[229] && f[320] && !f[461];
	assign leaf[4915] = f[693] && !f[229] && f[320] && f[461];
	assign leaf[4916] = f[693] && f[229] && !f[429];
	assign leaf[4917] = f[693] && f[229] && f[429] && !f[407];
	assign leaf[4918] = f[693] && f[229] && f[429] && f[407];
	
	// Tree 330, Classifier 0, Iteration: 33
	assign leaf[4919] = !f[571] && !f[436] && !f[360] && !f[512];
	assign leaf[4920] = !f[571] && !f[436] && !f[360] && f[512];
	assign leaf[4921] = !f[571] && !f[436] && f[360] && !f[275];
	assign leaf[4922] = !f[571] && !f[436] && f[360] && f[275];
	assign leaf[4923] = !f[571] && f[436] && !f[569] && !f[331];
	assign leaf[4924] = !f[571] && f[436] && !f[569] && f[331];
	assign leaf[4925] = !f[571] && f[436] && f[569] && !f[461];
	assign leaf[4926] = !f[571] && f[436] && f[569] && f[461];
	assign leaf[4927] = f[571] && !f[597] && !f[269] && !f[436];
	assign leaf[4928] = f[571] && !f[597] && !f[269] && f[436];
	assign leaf[4929] = f[571] && !f[597] && f[269] && !f[187];
	assign leaf[4930] = f[571] && !f[597] && f[269] && f[187];
	assign leaf[4931] = f[571] && f[597] && !f[608] && !f[300];
	assign leaf[4932] = f[571] && f[597] && !f[608] && f[300];
	assign leaf[4933] = f[571] && f[597] && f[608] && !f[498];
	assign leaf[4934] = f[571] && f[597] && f[608] && f[498];
	
	// Tree 331, Classifier 1, Iteration: 33
	assign leaf[4935] = !f[716] && !f[713] && !f[496] && !f[185];
	assign leaf[4936] = !f[716] && !f[713] && !f[496] && f[185];
	assign leaf[4937] = !f[716] && !f[713] && f[496] && !f[566];
	assign leaf[4938] = !f[716] && !f[713] && f[496] && f[566];
	assign leaf[4939] = !f[716] && f[713] && !f[345] && !f[407];
	assign leaf[4940] = !f[716] && f[713] && !f[345] && f[407];
	assign leaf[4941] = !f[716] && f[713] && f[345];
	assign leaf[4942] = f[716];
	
	// Tree 332, Classifier 2, Iteration: 33
	assign leaf[4943] = !f[713] && !f[710] && !f[95] && !f[322];
	assign leaf[4944] = !f[713] && !f[710] && !f[95] && f[322];
	assign leaf[4945] = !f[713] && !f[710] && f[95] && !f[262];
	assign leaf[4946] = !f[713] && !f[710] && f[95] && f[262];
	assign leaf[4947] = !f[713] && f[710];
	assign leaf[4948] = f[713] && !f[626];
	assign leaf[4949] = f[713] && f[626];
	
	// Tree 333, Classifier 3, Iteration: 33
	assign leaf[4950] = !f[712] && !f[535] && !f[657] && !f[458];
	assign leaf[4951] = !f[712] && !f[535] && !f[657] && f[458];
	assign leaf[4952] = !f[712] && !f[535] && f[657] && !f[709];
	assign leaf[4953] = !f[712] && !f[535] && f[657] && f[709];
	assign leaf[4954] = !f[712] && f[535] && !f[458] && !f[441];
	assign leaf[4955] = !f[712] && f[535] && !f[458] && f[441];
	assign leaf[4956] = !f[712] && f[535] && f[458] && !f[510];
	assign leaf[4957] = !f[712] && f[535] && f[458] && f[510];
	assign leaf[4958] = f[712] && !f[573] && !f[489] && !f[343];
	assign leaf[4959] = f[712] && !f[573] && !f[489] && f[343];
	assign leaf[4960] = f[712] && !f[573] && f[489] && !f[598];
	assign leaf[4961] = f[712] && !f[573] && f[489] && f[598];
	assign leaf[4962] = f[712] && f[573] && !f[488] && !f[429];
	assign leaf[4963] = f[712] && f[573] && !f[488] && f[429];
	assign leaf[4964] = f[712] && f[573] && f[488] && !f[599];
	assign leaf[4965] = f[712] && f[573] && f[488] && f[599];
	
	// Tree 334, Classifier 4, Iteration: 33
	assign leaf[4966] = !f[490] && !f[411] && !f[236] && !f[268];
	assign leaf[4967] = !f[490] && !f[411] && !f[236] && f[268];
	assign leaf[4968] = !f[490] && !f[411] && f[236] && !f[262];
	assign leaf[4969] = !f[490] && !f[411] && f[236] && f[262];
	assign leaf[4970] = !f[490] && f[411] && !f[323] && !f[397];
	assign leaf[4971] = !f[490] && f[411] && !f[323] && f[397];
	assign leaf[4972] = !f[490] && f[411] && f[323] && !f[435];
	assign leaf[4973] = !f[490] && f[411] && f[323] && f[435];
	assign leaf[4974] = f[490] && !f[348] && !f[346] && !f[344];
	assign leaf[4975] = f[490] && !f[348] && !f[346] && f[344];
	assign leaf[4976] = f[490] && !f[348] && f[346] && !f[243];
	assign leaf[4977] = f[490] && !f[348] && f[346] && f[243];
	assign leaf[4978] = f[490] && f[348] && !f[322] && !f[186];
	assign leaf[4979] = f[490] && f[348] && !f[322] && f[186];
	assign leaf[4980] = f[490] && f[348] && f[322] && !f[211];
	assign leaf[4981] = f[490] && f[348] && f[322] && f[211];
	
	// Tree 335, Classifier 5, Iteration: 33
	assign leaf[4982] = !f[434] && !f[464] && !f[713] && !f[120];
	assign leaf[4983] = !f[434] && !f[464] && !f[713] && f[120];
	assign leaf[4984] = !f[434] && !f[464] && f[713] && !f[465];
	assign leaf[4985] = !f[434] && !f[464] && f[713] && f[465];
	assign leaf[4986] = !f[434] && f[464] && !f[350] && !f[377];
	assign leaf[4987] = !f[434] && f[464] && !f[350] && f[377];
	assign leaf[4988] = !f[434] && f[464] && f[350] && !f[265];
	assign leaf[4989] = !f[434] && f[464] && f[350] && f[265];
	assign leaf[4990] = f[434] && !f[353] && !f[412] && !f[323];
	assign leaf[4991] = f[434] && !f[353] && !f[412] && f[323];
	assign leaf[4992] = f[434] && !f[353] && f[412] && !f[500];
	assign leaf[4993] = f[434] && !f[353] && f[412] && f[500];
	assign leaf[4994] = f[434] && f[353] && !f[347] && !f[304];
	assign leaf[4995] = f[434] && f[353] && !f[347] && f[304];
	assign leaf[4996] = f[434] && f[353] && f[347] && !f[276];
	assign leaf[4997] = f[434] && f[353] && f[347] && f[276];
	
	// Tree 336, Classifier 6, Iteration: 33
	assign leaf[4998] = !f[683] && !f[459] && !f[457] && !f[454];
	assign leaf[4999] = !f[683] && !f[459] && !f[457] && f[454];
	assign leaf[5000] = !f[683] && !f[459] && f[457] && !f[462];
	assign leaf[5001] = !f[683] && !f[459] && f[457] && f[462];
	assign leaf[5002] = !f[683] && f[459] && !f[375] && !f[292];
	assign leaf[5003] = !f[683] && f[459] && !f[375] && f[292];
	assign leaf[5004] = !f[683] && f[459] && f[375] && !f[303];
	assign leaf[5005] = !f[683] && f[459] && f[375] && f[303];
	assign leaf[5006] = f[683];
	
	// Tree 337, Classifier 7, Iteration: 33
	assign leaf[5007] = !f[242] && !f[411] && !f[177] && !f[231];
	assign leaf[5008] = !f[242] && !f[411] && !f[177] && f[231];
	assign leaf[5009] = !f[242] && !f[411] && f[177] && !f[492];
	assign leaf[5010] = !f[242] && !f[411] && f[177] && f[492];
	assign leaf[5011] = !f[242] && f[411] && !f[323] && !f[463];
	assign leaf[5012] = !f[242] && f[411] && !f[323] && f[463];
	assign leaf[5013] = !f[242] && f[411] && f[323] && !f[550];
	assign leaf[5014] = !f[242] && f[411] && f[323] && f[550];
	assign leaf[5015] = f[242] && !f[240] && !f[236] && !f[156];
	assign leaf[5016] = f[242] && !f[240] && !f[236] && f[156];
	assign leaf[5017] = f[242] && !f[240] && f[236] && !f[322];
	assign leaf[5018] = f[242] && !f[240] && f[236] && f[322];
	assign leaf[5019] = f[242] && f[240] && !f[349] && !f[325];
	assign leaf[5020] = f[242] && f[240] && !f[349] && f[325];
	assign leaf[5021] = f[242] && f[240] && f[349] && !f[267];
	assign leaf[5022] = f[242] && f[240] && f[349] && f[267];
	
	// Tree 338, Classifier 8, Iteration: 33
	assign leaf[5023] = !f[440] && !f[315] && !f[290] && !f[292];
	assign leaf[5024] = !f[440] && !f[315] && !f[290] && f[292];
	assign leaf[5025] = !f[440] && !f[315] && f[290] && !f[264];
	assign leaf[5026] = !f[440] && !f[315] && f[290] && f[264];
	assign leaf[5027] = !f[440] && f[315] && !f[489] && !f[288];
	assign leaf[5028] = !f[440] && f[315] && !f[489] && f[288];
	assign leaf[5029] = !f[440] && f[315] && f[489] && !f[634];
	assign leaf[5030] = !f[440] && f[315] && f[489] && f[634];
	assign leaf[5031] = f[440] && !f[576] && !f[567] && !f[514];
	assign leaf[5032] = f[440] && !f[576] && !f[567] && f[514];
	assign leaf[5033] = f[440] && !f[576] && f[567] && !f[681];
	assign leaf[5034] = f[440] && !f[576] && f[567] && f[681];
	assign leaf[5035] = f[440] && f[576] && !f[637] && !f[634];
	assign leaf[5036] = f[440] && f[576] && !f[637] && f[634];
	assign leaf[5037] = f[440] && f[576] && f[637] && !f[657];
	assign leaf[5038] = f[440] && f[576] && f[637] && f[657];
	
	// Tree 339, Classifier 9, Iteration: 33
	assign leaf[5039] = !f[436] && !f[465] && !f[667] && !f[492];
	assign leaf[5040] = !f[436] && !f[465] && !f[667] && f[492];
	assign leaf[5041] = !f[436] && !f[465] && f[667] && !f[454];
	assign leaf[5042] = !f[436] && !f[465] && f[667] && f[454];
	assign leaf[5043] = !f[436] && f[465] && !f[293] && !f[462];
	assign leaf[5044] = !f[436] && f[465] && !f[293] && f[462];
	assign leaf[5045] = !f[436] && f[465] && f[293] && !f[433];
	assign leaf[5046] = !f[436] && f[465] && f[293] && f[433];
	assign leaf[5047] = f[436] && !f[469] && !f[572] && !f[413];
	assign leaf[5048] = f[436] && !f[469] && !f[572] && f[413];
	assign leaf[5049] = f[436] && !f[469] && f[572] && !f[346];
	assign leaf[5050] = f[436] && !f[469] && f[572] && f[346];
	assign leaf[5051] = f[436] && f[469] && !f[357] && !f[692];
	assign leaf[5052] = f[436] && f[469] && !f[357] && f[692];
	assign leaf[5053] = f[436] && f[469] && f[357] && !f[347];
	assign leaf[5054] = f[436] && f[469] && f[357] && f[347];
	
	// Tree 340, Classifier 0, Iteration: 34
	assign leaf[5055] = !f[514] && !f[510] && !f[512] && !f[508];
	assign leaf[5056] = !f[514] && !f[510] && !f[512] && f[508];
	assign leaf[5057] = !f[514] && !f[510] && f[512] && !f[323];
	assign leaf[5058] = !f[514] && !f[510] && f[512] && f[323];
	assign leaf[5059] = !f[514] && f[510] && !f[246] && !f[272];
	assign leaf[5060] = !f[514] && f[510] && !f[246] && f[272];
	assign leaf[5061] = !f[514] && f[510] && f[246] && !f[379];
	assign leaf[5062] = !f[514] && f[510] && f[246] && f[379];
	assign leaf[5063] = f[514] && !f[656] && !f[359] && !f[520];
	assign leaf[5064] = f[514] && !f[656] && !f[359] && f[520];
	assign leaf[5065] = f[514] && !f[656] && f[359] && !f[398];
	assign leaf[5066] = f[514] && !f[656] && f[359] && f[398];
	assign leaf[5067] = f[514] && f[656] && !f[521] && !f[153];
	assign leaf[5068] = f[514] && f[656] && !f[521] && f[153];
	assign leaf[5069] = f[514] && f[656] && f[521] && !f[483];
	assign leaf[5070] = f[514] && f[656] && f[521] && f[483];
	
	// Tree 341, Classifier 1, Iteration: 34
	assign leaf[5071] = !f[537] && !f[407] && !f[463] && !f[548];
	assign leaf[5072] = !f[537] && !f[407] && !f[463] && f[548];
	assign leaf[5073] = !f[537] && !f[407] && f[463] && !f[460];
	assign leaf[5074] = !f[537] && !f[407] && f[463] && f[460];
	assign leaf[5075] = !f[537] && f[407] && !f[322] && !f[209];
	assign leaf[5076] = !f[537] && f[407] && !f[322] && f[209];
	assign leaf[5077] = !f[537] && f[407] && f[322] && !f[462];
	assign leaf[5078] = !f[537] && f[407] && f[322] && f[462];
	assign leaf[5079] = f[537] && !f[487];
	assign leaf[5080] = f[537] && f[487];
	
	// Tree 342, Classifier 2, Iteration: 34
	assign leaf[5081] = !f[639] && !f[677] && !f[351] && !f[372];
	assign leaf[5082] = !f[639] && !f[677] && !f[351] && f[372];
	assign leaf[5083] = !f[639] && !f[677] && f[351] && !f[487];
	assign leaf[5084] = !f[639] && !f[677] && f[351] && f[487];
	assign leaf[5085] = !f[639] && f[677] && !f[289];
	assign leaf[5086] = !f[639] && f[677] && f[289];
	assign leaf[5087] = f[639] && !f[554] && !f[371] && !f[569];
	assign leaf[5088] = f[639] && !f[554] && !f[371] && f[569];
	assign leaf[5089] = f[639] && !f[554] && f[371];
	assign leaf[5090] = f[639] && f[554] && !f[550] && !f[382];
	assign leaf[5091] = f[639] && f[554] && !f[550] && f[382];
	assign leaf[5092] = f[639] && f[554] && f[550];
	
	// Tree 343, Classifier 3, Iteration: 34
	assign leaf[5093] = !f[712] && !f[649] && !f[173] && !f[480];
	assign leaf[5094] = !f[712] && !f[649] && !f[173] && f[480];
	assign leaf[5095] = !f[712] && !f[649] && f[173] && !f[553];
	assign leaf[5096] = !f[712] && !f[649] && f[173] && f[553];
	assign leaf[5097] = !f[712] && f[649] && !f[539] && !f[320];
	assign leaf[5098] = !f[712] && f[649] && !f[539] && f[320];
	assign leaf[5099] = !f[712] && f[649] && f[539] && !f[375];
	assign leaf[5100] = !f[712] && f[649] && f[539] && f[375];
	assign leaf[5101] = f[712] && !f[600] && !f[489] && !f[519];
	assign leaf[5102] = f[712] && !f[600] && !f[489] && f[519];
	assign leaf[5103] = f[712] && !f[600] && f[489] && !f[403];
	assign leaf[5104] = f[712] && !f[600] && f[489] && f[403];
	assign leaf[5105] = f[712] && f[600] && !f[287] && !f[328];
	assign leaf[5106] = f[712] && f[600] && !f[287] && f[328];
	assign leaf[5107] = f[712] && f[600] && f[287];
	
	// Tree 344, Classifier 4, Iteration: 34
	assign leaf[5108] = !f[746] && !f[456] && !f[408] && !f[322];
	assign leaf[5109] = !f[746] && !f[456] && !f[408] && f[322];
	assign leaf[5110] = !f[746] && !f[456] && f[408] && !f[524];
	assign leaf[5111] = !f[746] && !f[456] && f[408] && f[524];
	assign leaf[5112] = !f[746] && f[456] && !f[439] && !f[494];
	assign leaf[5113] = !f[746] && f[456] && !f[439] && f[494];
	assign leaf[5114] = !f[746] && f[456] && f[439] && !f[513];
	assign leaf[5115] = !f[746] && f[456] && f[439] && f[513];
	assign leaf[5116] = f[746];
	
	// Tree 345, Classifier 5, Iteration: 34
	assign leaf[5117] = !f[228] && !f[191] && !f[248] && !f[269];
	assign leaf[5118] = !f[228] && !f[191] && !f[248] && f[269];
	assign leaf[5119] = !f[228] && !f[191] && f[248] && !f[269];
	assign leaf[5120] = !f[228] && !f[191] && f[248] && f[269];
	assign leaf[5121] = !f[228] && f[191] && !f[159] && !f[328];
	assign leaf[5122] = !f[228] && f[191] && !f[159] && f[328];
	assign leaf[5123] = !f[228] && f[191] && f[159] && !f[248];
	assign leaf[5124] = !f[228] && f[191] && f[159] && f[248];
	assign leaf[5125] = f[228] && !f[172];
	assign leaf[5126] = f[228] && f[172];
	
	// Tree 346, Classifier 6, Iteration: 34
	assign leaf[5127] = !f[683] && !f[234] && !f[151] && !f[326];
	assign leaf[5128] = !f[683] && !f[234] && !f[151] && f[326];
	assign leaf[5129] = !f[683] && !f[234] && f[151] && !f[398];
	assign leaf[5130] = !f[683] && !f[234] && f[151] && f[398];
	assign leaf[5131] = !f[683] && f[234] && !f[266] && !f[545];
	assign leaf[5132] = !f[683] && f[234] && !f[266] && f[545];
	assign leaf[5133] = !f[683] && f[234] && f[266] && !f[272];
	assign leaf[5134] = !f[683] && f[234] && f[266] && f[272];
	assign leaf[5135] = f[683];
	
	// Tree 347, Classifier 7, Iteration: 34
	assign leaf[5136] = !f[460] && !f[515] && !f[379] && !f[569];
	assign leaf[5137] = !f[460] && !f[515] && !f[379] && f[569];
	assign leaf[5138] = !f[460] && !f[515] && f[379] && !f[349];
	assign leaf[5139] = !f[460] && !f[515] && f[379] && f[349];
	assign leaf[5140] = !f[460] && f[515] && !f[678] && !f[234];
	assign leaf[5141] = !f[460] && f[515] && !f[678] && f[234];
	assign leaf[5142] = !f[460] && f[515] && f[678] && !f[262];
	assign leaf[5143] = !f[460] && f[515] && f[678] && f[262];
	assign leaf[5144] = f[460] && !f[372] && !f[374] && !f[342];
	assign leaf[5145] = f[460] && !f[372] && !f[374] && f[342];
	assign leaf[5146] = f[460] && !f[372] && f[374] && !f[497];
	assign leaf[5147] = f[460] && !f[372] && f[374] && f[497];
	assign leaf[5148] = f[460] && f[372] && !f[471] && !f[568];
	assign leaf[5149] = f[460] && f[372] && !f[471] && f[568];
	assign leaf[5150] = f[460] && f[372] && f[471] && !f[549];
	assign leaf[5151] = f[460] && f[372] && f[471] && f[549];
	
	// Tree 348, Classifier 8, Iteration: 34
	assign leaf[5152] = !f[248] && !f[350] && !f[517] && !f[514];
	assign leaf[5153] = !f[248] && !f[350] && !f[517] && f[514];
	assign leaf[5154] = !f[248] && !f[350] && f[517] && !f[456];
	assign leaf[5155] = !f[248] && !f[350] && f[517] && f[456];
	assign leaf[5156] = !f[248] && f[350] && !f[517] && !f[293];
	assign leaf[5157] = !f[248] && f[350] && !f[517] && f[293];
	assign leaf[5158] = !f[248] && f[350] && f[517] && !f[632];
	assign leaf[5159] = !f[248] && f[350] && f[517] && f[632];
	assign leaf[5160] = f[248] && !f[186] && !f[401] && !f[485];
	assign leaf[5161] = f[248] && !f[186] && !f[401] && f[485];
	assign leaf[5162] = f[248] && !f[186] && f[401] && !f[432];
	assign leaf[5163] = f[248] && !f[186] && f[401] && f[432];
	assign leaf[5164] = f[248] && f[186] && !f[577] && !f[181];
	assign leaf[5165] = f[248] && f[186] && !f[577] && f[181];
	assign leaf[5166] = f[248] && f[186] && f[577] && !f[328];
	assign leaf[5167] = f[248] && f[186] && f[577] && f[328];
	
	// Tree 349, Classifier 9, Iteration: 34
	assign leaf[5168] = !f[229] && !f[162] && !f[175] && !f[639];
	assign leaf[5169] = !f[229] && !f[162] && !f[175] && f[639];
	assign leaf[5170] = !f[229] && !f[162] && f[175] && !f[151];
	assign leaf[5171] = !f[229] && !f[162] && f[175] && f[151];
	assign leaf[5172] = !f[229] && f[162] && !f[679];
	assign leaf[5173] = !f[229] && f[162] && f[679];
	assign leaf[5174] = f[229] && !f[151] && !f[407] && !f[429];
	assign leaf[5175] = f[229] && !f[151] && !f[407] && f[429];
	assign leaf[5176] = f[229] && !f[151] && f[407];
	assign leaf[5177] = f[229] && f[151];
	
	// Tree 350, Classifier 0, Iteration: 35
	assign leaf[5178] = !f[240] && !f[377] && !f[436] && !f[321];
	assign leaf[5179] = !f[240] && !f[377] && !f[436] && f[321];
	assign leaf[5180] = !f[240] && !f[377] && f[436] && !f[270];
	assign leaf[5181] = !f[240] && !f[377] && f[436] && f[270];
	assign leaf[5182] = !f[240] && f[377] && !f[461] && !f[218];
	assign leaf[5183] = !f[240] && f[377] && !f[461] && f[218];
	assign leaf[5184] = !f[240] && f[377] && f[461] && !f[380];
	assign leaf[5185] = !f[240] && f[377] && f[461] && f[380];
	assign leaf[5186] = f[240] && !f[297] && !f[271] && !f[275];
	assign leaf[5187] = f[240] && !f[297] && !f[271] && f[275];
	assign leaf[5188] = f[240] && !f[297] && f[271] && !f[321];
	assign leaf[5189] = f[240] && !f[297] && f[271] && f[321];
	assign leaf[5190] = f[240] && f[297] && !f[486] && !f[606];
	assign leaf[5191] = f[240] && f[297] && !f[486] && f[606];
	assign leaf[5192] = f[240] && f[297] && f[486] && !f[375];
	assign leaf[5193] = f[240] && f[297] && f[486] && f[375];
	
	// Tree 351, Classifier 1, Iteration: 35
	assign leaf[5194] = !f[344] && !f[711] && !f[679] && !f[294];
	assign leaf[5195] = !f[344] && !f[711] && !f[679] && f[294];
	assign leaf[5196] = !f[344] && !f[711] && f[679] && !f[185];
	assign leaf[5197] = !f[344] && !f[711] && f[679] && f[185];
	assign leaf[5198] = !f[344] && f[711] && !f[710];
	assign leaf[5199] = !f[344] && f[711] && f[710];
	assign leaf[5200] = f[344] && !f[125] && !f[156];
	assign leaf[5201] = f[344] && !f[125] && f[156] && !f[293];
	assign leaf[5202] = f[344] && !f[125] && f[156] && f[293];
	assign leaf[5203] = f[344] && f[125];
	
	// Tree 352, Classifier 2, Iteration: 35
	assign leaf[5204] = !f[179] && !f[655] && !f[630] && !f[242];
	assign leaf[5205] = !f[179] && !f[655] && !f[630] && f[242];
	assign leaf[5206] = !f[179] && !f[655] && f[630] && !f[651];
	assign leaf[5207] = !f[179] && !f[655] && f[630] && f[651];
	assign leaf[5208] = !f[179] && f[655] && !f[606] && !f[596];
	assign leaf[5209] = !f[179] && f[655] && !f[606] && f[596];
	assign leaf[5210] = !f[179] && f[655] && f[606] && !f[601];
	assign leaf[5211] = !f[179] && f[655] && f[606] && f[601];
	assign leaf[5212] = f[179] && !f[599] && !f[341] && !f[666];
	assign leaf[5213] = f[179] && !f[599] && !f[341] && f[666];
	assign leaf[5214] = f[179] && !f[599] && f[341] && !f[583];
	assign leaf[5215] = f[179] && !f[599] && f[341] && f[583];
	assign leaf[5216] = f[179] && f[599] && !f[690] && !f[409];
	assign leaf[5217] = f[179] && f[599] && !f[690] && f[409];
	assign leaf[5218] = f[179] && f[599] && f[690] && !f[636];
	assign leaf[5219] = f[179] && f[599] && f[690] && f[636];
	
	// Tree 353, Classifier 3, Iteration: 35
	assign leaf[5220] = !f[373] && !f[523] && !f[320] && !f[327];
	assign leaf[5221] = !f[373] && !f[523] && !f[320] && f[327];
	assign leaf[5222] = !f[373] && !f[523] && f[320] && !f[126];
	assign leaf[5223] = !f[373] && !f[523] && f[320] && f[126];
	assign leaf[5224] = !f[373] && f[523] && !f[238] && !f[263];
	assign leaf[5225] = !f[373] && f[523] && !f[238] && f[263];
	assign leaf[5226] = !f[373] && f[523] && f[238] && !f[161];
	assign leaf[5227] = !f[373] && f[523] && f[238] && f[161];
	assign leaf[5228] = f[373] && !f[288] && !f[526] && !f[154];
	assign leaf[5229] = f[373] && !f[288] && !f[526] && f[154];
	assign leaf[5230] = f[373] && !f[288] && f[526] && !f[293];
	assign leaf[5231] = f[373] && !f[288] && f[526] && f[293];
	assign leaf[5232] = f[373] && f[288] && !f[264] && !f[316];
	assign leaf[5233] = f[373] && f[288] && !f[264] && f[316];
	assign leaf[5234] = f[373] && f[288] && f[264] && !f[469];
	assign leaf[5235] = f[373] && f[288] && f[264] && f[469];
	
	// Tree 354, Classifier 4, Iteration: 35
	assign leaf[5236] = !f[740] && !f[185] && !f[183] && !f[294];
	assign leaf[5237] = !f[740] && !f[185] && !f[183] && f[294];
	assign leaf[5238] = !f[740] && !f[185] && f[183] && !f[180];
	assign leaf[5239] = !f[740] && !f[185] && f[183] && f[180];
	assign leaf[5240] = !f[740] && f[185] && !f[296] && !f[294];
	assign leaf[5241] = !f[740] && f[185] && !f[296] && f[294];
	assign leaf[5242] = !f[740] && f[185] && f[296] && !f[182];
	assign leaf[5243] = !f[740] && f[185] && f[296] && f[182];
	assign leaf[5244] = f[740] && !f[240];
	assign leaf[5245] = f[740] && f[240];
	
	// Tree 355, Classifier 5, Iteration: 35
	assign leaf[5246] = !f[188] && !f[245] && !f[240] && !f[157];
	assign leaf[5247] = !f[188] && !f[245] && !f[240] && f[157];
	assign leaf[5248] = !f[188] && !f[245] && f[240] && !f[236];
	assign leaf[5249] = !f[188] && !f[245] && f[240] && f[236];
	assign leaf[5250] = !f[188] && f[245] && !f[328] && !f[359];
	assign leaf[5251] = !f[188] && f[245] && !f[328] && f[359];
	assign leaf[5252] = !f[188] && f[245] && f[328] && !f[276];
	assign leaf[5253] = !f[188] && f[245] && f[328] && f[276];
	assign leaf[5254] = f[188] && !f[213] && !f[216] && !f[246];
	assign leaf[5255] = f[188] && !f[213] && !f[216] && f[246];
	assign leaf[5256] = f[188] && !f[213] && f[216] && !f[192];
	assign leaf[5257] = f[188] && !f[213] && f[216] && f[192];
	assign leaf[5258] = f[188] && f[213] && !f[300] && !f[303];
	assign leaf[5259] = f[188] && f[213] && !f[300] && f[303];
	assign leaf[5260] = f[188] && f[213] && f[300] && !f[688];
	assign leaf[5261] = f[188] && f[213] && f[300] && f[688];
	
	// Tree 356, Classifier 6, Iteration: 35
	assign leaf[5262] = !f[601] && !f[64] && !f[295] && !f[241];
	assign leaf[5263] = !f[601] && !f[64] && !f[295] && f[241];
	assign leaf[5264] = !f[601] && !f[64] && f[295] && !f[132];
	assign leaf[5265] = !f[601] && !f[64] && f[295] && f[132];
	assign leaf[5266] = !f[601] && f[64];
	assign leaf[5267] = f[601] && !f[486] && !f[455] && !f[516];
	assign leaf[5268] = f[601] && !f[486] && !f[455] && f[516];
	assign leaf[5269] = f[601] && !f[486] && f[455] && !f[370];
	assign leaf[5270] = f[601] && !f[486] && f[455] && f[370];
	assign leaf[5271] = f[601] && f[486] && !f[374] && !f[181];
	assign leaf[5272] = f[601] && f[486] && !f[374] && f[181];
	assign leaf[5273] = f[601] && f[486] && f[374] && !f[458];
	assign leaf[5274] = f[601] && f[486] && f[374] && f[458];
	
	// Tree 357, Classifier 7, Iteration: 35
	assign leaf[5275] = !f[555] && !f[129] && !f[635] && !f[437];
	assign leaf[5276] = !f[555] && !f[129] && !f[635] && f[437];
	assign leaf[5277] = !f[555] && !f[129] && f[635] && !f[319];
	assign leaf[5278] = !f[555] && !f[129] && f[635] && f[319];
	assign leaf[5279] = !f[555] && f[129];
	assign leaf[5280] = f[555] && !f[540];
	assign leaf[5281] = f[555] && f[540];
	
	// Tree 358, Classifier 8, Iteration: 35
	assign leaf[5282] = !f[248] && !f[156] && !f[542] && !f[544];
	assign leaf[5283] = !f[248] && !f[156] && !f[542] && f[544];
	assign leaf[5284] = !f[248] && !f[156] && f[542] && !f[455];
	assign leaf[5285] = !f[248] && !f[156] && f[542] && f[455];
	assign leaf[5286] = !f[248] && f[156] && !f[212] && !f[266];
	assign leaf[5287] = !f[248] && f[156] && !f[212] && f[266];
	assign leaf[5288] = !f[248] && f[156] && f[212] && !f[576];
	assign leaf[5289] = !f[248] && f[156] && f[212] && f[576];
	assign leaf[5290] = f[248] && !f[347] && !f[322] && !f[575];
	assign leaf[5291] = f[248] && !f[347] && !f[322] && f[575];
	assign leaf[5292] = f[248] && !f[347] && f[322] && !f[352];
	assign leaf[5293] = f[248] && !f[347] && f[322] && f[352];
	assign leaf[5294] = f[248] && f[347] && !f[383] && !f[374];
	assign leaf[5295] = f[248] && f[347] && !f[383] && f[374];
	assign leaf[5296] = f[248] && f[347] && f[383] && !f[371];
	assign leaf[5297] = f[248] && f[347] && f[383] && f[371];
	
	// Tree 359, Classifier 9, Iteration: 35
	assign leaf[5298] = !f[742] && !f[632] && !f[688] && !f[542];
	assign leaf[5299] = !f[742] && !f[632] && !f[688] && f[542];
	assign leaf[5300] = !f[742] && !f[632] && f[688] && !f[662];
	assign leaf[5301] = !f[742] && !f[632] && f[688] && f[662];
	assign leaf[5302] = !f[742] && f[632] && !f[493] && !f[517];
	assign leaf[5303] = !f[742] && f[632] && !f[493] && f[517];
	assign leaf[5304] = !f[742] && f[632] && f[493] && !f[182];
	assign leaf[5305] = !f[742] && f[632] && f[493] && f[182];
	assign leaf[5306] = f[742] && !f[634] && !f[204] && !f[290];
	assign leaf[5307] = f[742] && !f[634] && !f[204] && f[290];
	assign leaf[5308] = f[742] && !f[634] && f[204];
	assign leaf[5309] = f[742] && f[634];
	
	// Tree 360, Classifier 0, Iteration: 36
	assign leaf[5310] = !f[711] && !f[609] && !f[177] && !f[415];
	assign leaf[5311] = !f[711] && !f[609] && !f[177] && f[415];
	assign leaf[5312] = !f[711] && !f[609] && f[177] && !f[572];
	assign leaf[5313] = !f[711] && !f[609] && f[177] && f[572];
	assign leaf[5314] = !f[711] && f[609] && !f[471] && !f[662];
	assign leaf[5315] = !f[711] && f[609] && !f[471] && f[662];
	assign leaf[5316] = !f[711] && f[609] && f[471] && !f[346];
	assign leaf[5317] = !f[711] && f[609] && f[471] && f[346];
	assign leaf[5318] = f[711] && !f[573];
	assign leaf[5319] = f[711] && f[573];
	
	// Tree 361, Classifier 1, Iteration: 36
	assign leaf[5320] = !f[440] && !f[710] && !f[407] && !f[463];
	assign leaf[5321] = !f[440] && !f[710] && !f[407] && f[463];
	assign leaf[5322] = !f[440] && !f[710] && f[407] && !f[578];
	assign leaf[5323] = !f[440] && !f[710] && f[407] && f[578];
	assign leaf[5324] = !f[440] && f[710] && !f[238];
	assign leaf[5325] = !f[440] && f[710] && f[238];
	assign leaf[5326] = f[440];
	
	// Tree 362, Classifier 2, Iteration: 36
	assign leaf[5327] = !f[397] && !f[388] && !f[374] && !f[349];
	assign leaf[5328] = !f[397] && !f[388] && !f[374] && f[349];
	assign leaf[5329] = !f[397] && !f[388] && f[374] && !f[318];
	assign leaf[5330] = !f[397] && !f[388] && f[374] && f[318];
	assign leaf[5331] = !f[397] && f[388] && !f[399] && !f[214];
	assign leaf[5332] = !f[397] && f[388] && !f[399] && f[214];
	assign leaf[5333] = !f[397] && f[388] && f[399] && !f[343];
	assign leaf[5334] = !f[397] && f[388] && f[399] && f[343];
	assign leaf[5335] = f[397] && !f[374] && !f[426] && !f[495];
	assign leaf[5336] = f[397] && !f[374] && !f[426] && f[495];
	assign leaf[5337] = f[397] && !f[374] && f[426] && !f[508];
	assign leaf[5338] = f[397] && !f[374] && f[426] && f[508];
	assign leaf[5339] = f[397] && f[374] && !f[287] && !f[521];
	assign leaf[5340] = f[397] && f[374] && !f[287] && f[521];
	assign leaf[5341] = f[397] && f[374] && f[287];
	
	// Tree 363, Classifier 3, Iteration: 36
	assign leaf[5342] = !f[386] && !f[269] && !f[129] && !f[491];
	assign leaf[5343] = !f[386] && !f[269] && !f[129] && f[491];
	assign leaf[5344] = !f[386] && !f[269] && f[129] && !f[272];
	assign leaf[5345] = !f[386] && !f[269] && f[129] && f[272];
	assign leaf[5346] = !f[386] && f[269] && !f[99] && !f[572];
	assign leaf[5347] = !f[386] && f[269] && !f[99] && f[572];
	assign leaf[5348] = !f[386] && f[269] && f[99] && !f[179];
	assign leaf[5349] = !f[386] && f[269] && f[99] && f[179];
	assign leaf[5350] = f[386] && !f[354];
	assign leaf[5351] = f[386] && f[354] && !f[149] && !f[381];
	assign leaf[5352] = f[386] && f[354] && !f[149] && f[381];
	assign leaf[5353] = f[386] && f[354] && f[149] && !f[267];
	assign leaf[5354] = f[386] && f[354] && f[149] && f[267];
	
	// Tree 364, Classifier 4, Iteration: 36
	assign leaf[5355] = !f[744] && !f[128] && !f[739] && !f[747];
	assign leaf[5356] = !f[744] && !f[128] && !f[739] && f[747];
	assign leaf[5357] = !f[744] && !f[128] && f[739] && !f[412];
	assign leaf[5358] = !f[744] && !f[128] && f[739] && f[412];
	assign leaf[5359] = !f[744] && f[128] && !f[239] && !f[433];
	assign leaf[5360] = !f[744] && f[128] && !f[239] && f[433];
	assign leaf[5361] = !f[744] && f[128] && f[239] && !f[628];
	assign leaf[5362] = !f[744] && f[128] && f[239] && f[628];
	assign leaf[5363] = f[744] && !f[455] && !f[411];
	assign leaf[5364] = f[744] && !f[455] && f[411];
	assign leaf[5365] = f[744] && f[455];
	
	// Tree 365, Classifier 5, Iteration: 36
	assign leaf[5366] = !f[102] && !f[565] && !f[289] && !f[481];
	assign leaf[5367] = !f[102] && !f[565] && !f[289] && f[481];
	assign leaf[5368] = !f[102] && !f[565] && f[289] && !f[178];
	assign leaf[5369] = !f[102] && !f[565] && f[289] && f[178];
	assign leaf[5370] = !f[102] && f[565] && !f[302] && !f[267];
	assign leaf[5371] = !f[102] && f[565] && !f[302] && f[267];
	assign leaf[5372] = !f[102] && f[565] && f[302] && !f[271];
	assign leaf[5373] = !f[102] && f[565] && f[302] && f[271];
	assign leaf[5374] = f[102] && !f[242] && !f[324] && !f[206];
	assign leaf[5375] = f[102] && !f[242] && !f[324] && f[206];
	assign leaf[5376] = f[102] && !f[242] && f[324] && !f[291];
	assign leaf[5377] = f[102] && !f[242] && f[324] && f[291];
	assign leaf[5378] = f[102] && f[242] && !f[347];
	assign leaf[5379] = f[102] && f[242] && f[347];
	
	// Tree 366, Classifier 6, Iteration: 36
	assign leaf[5380] = !f[637] && !f[299] && !f[301] && !f[324];
	assign leaf[5381] = !f[637] && !f[299] && !f[301] && f[324];
	assign leaf[5382] = !f[637] && !f[299] && f[301] && !f[122];
	assign leaf[5383] = !f[637] && !f[299] && f[301] && f[122];
	assign leaf[5384] = !f[637] && f[299] && !f[382] && !f[176];
	assign leaf[5385] = !f[637] && f[299] && !f[382] && f[176];
	assign leaf[5386] = !f[637] && f[299] && f[382] && !f[357];
	assign leaf[5387] = !f[637] && f[299] && f[382] && f[357];
	assign leaf[5388] = f[637] && !f[511] && !f[526] && !f[125];
	assign leaf[5389] = f[637] && !f[511] && !f[526] && f[125];
	assign leaf[5390] = f[637] && !f[511] && f[526];
	assign leaf[5391] = f[637] && f[511] && !f[263];
	assign leaf[5392] = f[637] && f[511] && f[263];
	
	// Tree 367, Classifier 7, Iteration: 36
	assign leaf[5393] = !f[127] && !f[677] && !f[595] && !f[515];
	assign leaf[5394] = !f[127] && !f[677] && !f[595] && f[515];
	assign leaf[5395] = !f[127] && !f[677] && f[595] && !f[406];
	assign leaf[5396] = !f[127] && !f[677] && f[595] && f[406];
	assign leaf[5397] = !f[127] && f[677] && !f[576] && !f[541];
	assign leaf[5398] = !f[127] && f[677] && !f[576] && f[541];
	assign leaf[5399] = !f[127] && f[677] && f[576];
	assign leaf[5400] = f[127] && !f[539];
	assign leaf[5401] = f[127] && f[539];
	
	// Tree 368, Classifier 8, Iteration: 36
	assign leaf[5402] = !f[340] && !f[399] && !f[317] && !f[291];
	assign leaf[5403] = !f[340] && !f[399] && !f[317] && f[291];
	assign leaf[5404] = !f[340] && !f[399] && f[317] && !f[403];
	assign leaf[5405] = !f[340] && !f[399] && f[317] && f[403];
	assign leaf[5406] = !f[340] && f[399] && !f[493] && !f[510];
	assign leaf[5407] = !f[340] && f[399] && !f[493] && f[510];
	assign leaf[5408] = !f[340] && f[399] && f[493] && !f[346];
	assign leaf[5409] = !f[340] && f[399] && f[493] && f[346];
	assign leaf[5410] = f[340] && !f[464];
	assign leaf[5411] = f[340] && f[464] && !f[152] && !f[546];
	assign leaf[5412] = f[340] && f[464] && !f[152] && f[546];
	assign leaf[5413] = f[340] && f[464] && f[152];
	
	// Tree 369, Classifier 9, Iteration: 36
	assign leaf[5414] = !f[356] && !f[468] && !f[412] && !f[244];
	assign leaf[5415] = !f[356] && !f[468] && !f[412] && f[244];
	assign leaf[5416] = !f[356] && !f[468] && f[412] && !f[495];
	assign leaf[5417] = !f[356] && !f[468] && f[412] && f[495];
	assign leaf[5418] = !f[356] && f[468] && !f[408] && !f[287];
	assign leaf[5419] = !f[356] && f[468] && !f[408] && f[287];
	assign leaf[5420] = !f[356] && f[468] && f[408] && !f[694];
	assign leaf[5421] = !f[356] && f[468] && f[408] && f[694];
	assign leaf[5422] = f[356] && !f[411] && !f[741] && !f[437];
	assign leaf[5423] = f[356] && !f[411] && !f[741] && f[437];
	assign leaf[5424] = f[356] && !f[411] && f[741];
	assign leaf[5425] = f[356] && f[411] && !f[213] && !f[185];
	assign leaf[5426] = f[356] && f[411] && !f[213] && f[185];
	assign leaf[5427] = f[356] && f[411] && f[213] && !f[295];
	assign leaf[5428] = f[356] && f[411] && f[213] && f[295];
	
	// Tree 370, Classifier 0, Iteration: 37
	assign leaf[5429] = !f[213] && !f[408] && !f[377] && !f[461];
	assign leaf[5430] = !f[213] && !f[408] && !f[377] && f[461];
	assign leaf[5431] = !f[213] && !f[408] && f[377] && !f[437];
	assign leaf[5432] = !f[213] && !f[408] && f[377] && f[437];
	assign leaf[5433] = !f[213] && f[408] && !f[268] && !f[151];
	assign leaf[5434] = !f[213] && f[408] && !f[268] && f[151];
	assign leaf[5435] = !f[213] && f[408] && f[268] && !f[490];
	assign leaf[5436] = !f[213] && f[408] && f[268] && f[490];
	assign leaf[5437] = f[213] && !f[711] && !f[634] && !f[580];
	assign leaf[5438] = f[213] && !f[711] && !f[634] && f[580];
	assign leaf[5439] = f[213] && !f[711] && f[634] && !f[466];
	assign leaf[5440] = f[213] && !f[711] && f[634] && f[466];
	assign leaf[5441] = f[213] && f[711] && !f[295];
	assign leaf[5442] = f[213] && f[711] && f[295];
	
	// Tree 371, Classifier 1, Iteration: 37
	assign leaf[5443] = !f[511] && !f[713] && !f[537] && !f[316];
	assign leaf[5444] = !f[511] && !f[713] && !f[537] && f[316];
	assign leaf[5445] = !f[511] && !f[713] && f[537];
	assign leaf[5446] = !f[511] && f[713] && !f[659] && !f[186];
	assign leaf[5447] = !f[511] && f[713] && !f[659] && f[186];
	assign leaf[5448] = !f[511] && f[713] && f[659] && !f[404];
	assign leaf[5449] = !f[511] && f[713] && f[659] && f[404];
	assign leaf[5450] = f[511] && !f[430] && !f[549] && !f[408];
	assign leaf[5451] = f[511] && !f[430] && !f[549] && f[408];
	assign leaf[5452] = f[511] && !f[430] && f[549];
	assign leaf[5453] = f[511] && f[430] && !f[242];
	assign leaf[5454] = f[511] && f[430] && f[242] && !f[600];
	assign leaf[5455] = f[511] && f[430] && f[242] && f[600];
	
	// Tree 372, Classifier 2, Iteration: 37
	assign leaf[5456] = !f[473] && !f[293] && !f[289] && !f[427];
	assign leaf[5457] = !f[473] && !f[293] && !f[289] && f[427];
	assign leaf[5458] = !f[473] && !f[293] && f[289] && !f[373];
	assign leaf[5459] = !f[473] && !f[293] && f[289] && f[373];
	assign leaf[5460] = !f[473] && f[293] && !f[388] && !f[620];
	assign leaf[5461] = !f[473] && f[293] && !f[388] && f[620];
	assign leaf[5462] = !f[473] && f[293] && f[388] && !f[359];
	assign leaf[5463] = !f[473] && f[293] && f[388] && f[359];
	assign leaf[5464] = f[473] && !f[416] && !f[485];
	assign leaf[5465] = f[473] && !f[416] && f[485] && !f[400];
	assign leaf[5466] = f[473] && !f[416] && f[485] && f[400];
	assign leaf[5467] = f[473] && f[416];
	
	// Tree 373, Classifier 3, Iteration: 37
	assign leaf[5468] = !f[708] && !f[550] && !f[553] && !f[98];
	assign leaf[5469] = !f[708] && !f[550] && !f[553] && f[98];
	assign leaf[5470] = !f[708] && !f[550] && f[553] && !f[547];
	assign leaf[5471] = !f[708] && !f[550] && f[553] && f[547];
	assign leaf[5472] = !f[708] && f[550] && !f[401] && !f[544];
	assign leaf[5473] = !f[708] && f[550] && !f[401] && f[544];
	assign leaf[5474] = !f[708] && f[550] && f[401] && !f[455];
	assign leaf[5475] = !f[708] && f[550] && f[401] && f[455];
	assign leaf[5476] = f[708] && !f[576] && !f[599] && !f[293];
	assign leaf[5477] = f[708] && !f[576] && !f[599] && f[293];
	assign leaf[5478] = f[708] && !f[576] && f[599] && !f[516];
	assign leaf[5479] = f[708] && !f[576] && f[599] && f[516];
	assign leaf[5480] = f[708] && f[576] && !f[376];
	assign leaf[5481] = f[708] && f[576] && f[376] && !f[380];
	assign leaf[5482] = f[708] && f[576] && f[376] && f[380];
	
	// Tree 374, Classifier 4, Iteration: 37
	assign leaf[5483] = !f[737] && !f[743] && !f[180] && !f[236];
	assign leaf[5484] = !f[737] && !f[743] && !f[180] && f[236];
	assign leaf[5485] = !f[737] && !f[743] && f[180] && !f[183];
	assign leaf[5486] = !f[737] && !f[743] && f[180] && f[183];
	assign leaf[5487] = !f[737] && f[743] && !f[298] && !f[353];
	assign leaf[5488] = !f[737] && f[743] && !f[298] && f[353];
	assign leaf[5489] = !f[737] && f[743] && f[298] && !f[490];
	assign leaf[5490] = !f[737] && f[743] && f[298] && f[490];
	assign leaf[5491] = f[737] && !f[385];
	assign leaf[5492] = f[737] && f[385];
	
	// Tree 375, Classifier 5, Iteration: 37
	assign leaf[5493] = !f[333] && !f[485] && !f[160] && !f[218];
	assign leaf[5494] = !f[333] && !f[485] && !f[160] && f[218];
	assign leaf[5495] = !f[333] && !f[485] && f[160] && !f[243];
	assign leaf[5496] = !f[333] && !f[485] && f[160] && f[243];
	assign leaf[5497] = !f[333] && f[485] && !f[158] && !f[244];
	assign leaf[5498] = !f[333] && f[485] && !f[158] && f[244];
	assign leaf[5499] = !f[333] && f[485] && f[158] && !f[577];
	assign leaf[5500] = !f[333] && f[485] && f[158] && f[577];
	assign leaf[5501] = f[333] && !f[330];
	assign leaf[5502] = f[333] && f[330] && !f[571];
	assign leaf[5503] = f[333] && f[330] && f[571];
	
	// Tree 376, Classifier 6, Iteration: 37
	assign leaf[5504] = !f[653] && !f[689] && !f[517] && !f[151];
	assign leaf[5505] = !f[653] && !f[689] && !f[517] && f[151];
	assign leaf[5506] = !f[653] && !f[689] && f[517] && !f[240];
	assign leaf[5507] = !f[653] && !f[689] && f[517] && f[240];
	assign leaf[5508] = !f[653] && f[689] && !f[598];
	assign leaf[5509] = !f[653] && f[689] && f[598];
	assign leaf[5510] = f[653] && !f[162] && !f[627] && !f[519];
	assign leaf[5511] = f[653] && !f[162] && !f[627] && f[519];
	assign leaf[5512] = f[653] && !f[162] && f[627];
	assign leaf[5513] = f[653] && f[162] && !f[490] && !f[539];
	assign leaf[5514] = f[653] && f[162] && !f[490] && f[539];
	assign leaf[5515] = f[653] && f[162] && f[490];
	
	// Tree 377, Classifier 7, Iteration: 37
	assign leaf[5516] = !f[256] && !f[663] && !f[349] && !f[433];
	assign leaf[5517] = !f[256] && !f[663] && !f[349] && f[433];
	assign leaf[5518] = !f[256] && !f[663] && f[349] && !f[384];
	assign leaf[5519] = !f[256] && !f[663] && f[349] && f[384];
	assign leaf[5520] = !f[256] && f[663] && !f[263] && !f[178];
	assign leaf[5521] = !f[256] && f[663] && !f[263] && f[178];
	assign leaf[5522] = !f[256] && f[663] && f[263] && !f[489];
	assign leaf[5523] = !f[256] && f[663] && f[263] && f[489];
	assign leaf[5524] = f[256] && !f[287] && !f[659] && !f[494];
	assign leaf[5525] = f[256] && !f[287] && !f[659] && f[494];
	assign leaf[5526] = f[256] && !f[287] && f[659];
	assign leaf[5527] = f[256] && f[287] && !f[554] && !f[294];
	assign leaf[5528] = f[256] && f[287] && !f[554] && f[294];
	assign leaf[5529] = f[256] && f[287] && f[554];
	
	// Tree 378, Classifier 8, Iteration: 37
	assign leaf[5530] = !f[679] && !f[273] && !f[710] && !f[438];
	assign leaf[5531] = !f[679] && !f[273] && !f[710] && f[438];
	assign leaf[5532] = !f[679] && !f[273] && f[710] && !f[542];
	assign leaf[5533] = !f[679] && !f[273] && f[710] && f[542];
	assign leaf[5534] = !f[679] && f[273] && !f[480] && !f[243];
	assign leaf[5535] = !f[679] && f[273] && !f[480] && f[243];
	assign leaf[5536] = !f[679] && f[273] && f[480] && !f[633];
	assign leaf[5537] = !f[679] && f[273] && f[480] && f[633];
	assign leaf[5538] = f[679] && !f[540] && !f[711] && !f[538];
	assign leaf[5539] = f[679] && !f[540] && !f[711] && f[538];
	assign leaf[5540] = f[679] && !f[540] && f[711] && !f[182];
	assign leaf[5541] = f[679] && !f[540] && f[711] && f[182];
	assign leaf[5542] = f[679] && f[540] && !f[681] && !f[621];
	assign leaf[5543] = f[679] && f[540] && !f[681] && f[621];
	assign leaf[5544] = f[679] && f[540] && f[681] && !f[232];
	assign leaf[5545] = f[679] && f[540] && f[681] && f[232];
	
	// Tree 379, Classifier 9, Iteration: 37
	assign leaf[5546] = !f[191] && !f[319] && !f[371] && !f[345];
	assign leaf[5547] = !f[191] && !f[319] && !f[371] && f[345];
	assign leaf[5548] = !f[191] && !f[319] && f[371] && !f[345];
	assign leaf[5549] = !f[191] && !f[319] && f[371] && f[345];
	assign leaf[5550] = !f[191] && f[319] && !f[522] && !f[467];
	assign leaf[5551] = !f[191] && f[319] && !f[522] && f[467];
	assign leaf[5552] = !f[191] && f[319] && f[522] && !f[410];
	assign leaf[5553] = !f[191] && f[319] && f[522] && f[410];
	assign leaf[5554] = f[191] && !f[273] && !f[399];
	assign leaf[5555] = f[191] && !f[273] && f[399];
	assign leaf[5556] = f[191] && f[273] && !f[482];
	assign leaf[5557] = f[191] && f[273] && f[482];
	
	// Tree 380, Classifier 0, Iteration: 38
	assign leaf[5558] = !f[378] && !f[517] && !f[629] && !f[684];
	assign leaf[5559] = !f[378] && !f[517] && !f[629] && f[684];
	assign leaf[5560] = !f[378] && !f[517] && f[629] && !f[323];
	assign leaf[5561] = !f[378] && !f[517] && f[629] && f[323];
	assign leaf[5562] = !f[378] && f[517] && !f[427] && !f[377];
	assign leaf[5563] = !f[378] && f[517] && !f[427] && f[377];
	assign leaf[5564] = !f[378] && f[517] && f[427] && !f[330];
	assign leaf[5565] = !f[378] && f[517] && f[427] && f[330];
	assign leaf[5566] = f[378] && !f[216] && !f[376] && !f[606];
	assign leaf[5567] = f[378] && !f[216] && !f[376] && f[606];
	assign leaf[5568] = f[378] && !f[216] && f[376] && !f[406];
	assign leaf[5569] = f[378] && !f[216] && f[376] && f[406];
	assign leaf[5570] = f[378] && f[216] && !f[568] && !f[570];
	assign leaf[5571] = f[378] && f[216] && !f[568] && f[570];
	assign leaf[5572] = f[378] && f[216] && f[568] && !f[326];
	assign leaf[5573] = f[378] && f[216] && f[568] && f[326];
	
	// Tree 381, Classifier 1, Iteration: 38
	assign leaf[5574] = !f[621] && !f[204] && !f[565] && !f[628];
	assign leaf[5575] = !f[621] && !f[204] && !f[565] && f[628];
	assign leaf[5576] = !f[621] && !f[204] && f[565] && !f[488];
	assign leaf[5577] = !f[621] && !f[204] && f[565] && f[488];
	assign leaf[5578] = !f[621] && f[204] && !f[625] && !f[291];
	assign leaf[5579] = !f[621] && f[204] && !f[625] && f[291];
	assign leaf[5580] = !f[621] && f[204] && f[625] && !f[150];
	assign leaf[5581] = !f[621] && f[204] && f[625] && f[150];
	assign leaf[5582] = f[621] && !f[605] && !f[600] && !f[219];
	assign leaf[5583] = f[621] && !f[605] && !f[600] && f[219];
	assign leaf[5584] = f[621] && !f[605] && f[600];
	assign leaf[5585] = f[621] && f[605];
	
	// Tree 382, Classifier 2, Iteration: 38
	assign leaf[5586] = !f[324] && !f[485] && !f[298] && !f[380];
	assign leaf[5587] = !f[324] && !f[485] && !f[298] && f[380];
	assign leaf[5588] = !f[324] && !f[485] && f[298] && !f[432];
	assign leaf[5589] = !f[324] && !f[485] && f[298] && f[432];
	assign leaf[5590] = !f[324] && f[485] && !f[285] && !f[343];
	assign leaf[5591] = !f[324] && f[485] && !f[285] && f[343];
	assign leaf[5592] = !f[324] && f[485] && f[285] && !f[231];
	assign leaf[5593] = !f[324] && f[485] && f[285] && f[231];
	assign leaf[5594] = f[324] && !f[411] && !f[271] && !f[159];
	assign leaf[5595] = f[324] && !f[411] && !f[271] && f[159];
	assign leaf[5596] = f[324] && !f[411] && f[271] && !f[606];
	assign leaf[5597] = f[324] && !f[411] && f[271] && f[606];
	assign leaf[5598] = f[324] && f[411] && !f[415] && !f[172];
	assign leaf[5599] = f[324] && f[411] && !f[415] && f[172];
	assign leaf[5600] = f[324] && f[411] && f[415] && !f[243];
	assign leaf[5601] = f[324] && f[411] && f[415] && f[243];
	
	// Tree 383, Classifier 3, Iteration: 38
	assign leaf[5602] = !f[457] && !f[96] && !f[406] && !f[461];
	assign leaf[5603] = !f[457] && !f[96] && !f[406] && f[461];
	assign leaf[5604] = !f[457] && !f[96] && f[406] && !f[300];
	assign leaf[5605] = !f[457] && !f[96] && f[406] && f[300];
	assign leaf[5606] = !f[457] && f[96] && !f[265] && !f[568];
	assign leaf[5607] = !f[457] && f[96] && !f[265] && f[568];
	assign leaf[5608] = !f[457] && f[96] && f[265] && !f[180];
	assign leaf[5609] = !f[457] && f[96] && f[265] && f[180];
	assign leaf[5610] = f[457] && !f[235] && !f[578] && !f[508];
	assign leaf[5611] = f[457] && !f[235] && !f[578] && f[508];
	assign leaf[5612] = f[457] && !f[235] && f[578] && !f[324];
	assign leaf[5613] = f[457] && !f[235] && f[578] && f[324];
	assign leaf[5614] = f[457] && f[235] && !f[406] && !f[598];
	assign leaf[5615] = f[457] && f[235] && !f[406] && f[598];
	assign leaf[5616] = f[457] && f[235] && f[406] && !f[346];
	assign leaf[5617] = f[457] && f[235] && f[406] && f[346];
	
	// Tree 384, Classifier 4, Iteration: 38
	assign leaf[5618] = !f[332] && !f[737] && !f[185] && !f[187];
	assign leaf[5619] = !f[332] && !f[737] && !f[185] && f[187];
	assign leaf[5620] = !f[332] && !f[737] && f[185] && !f[182];
	assign leaf[5621] = !f[332] && !f[737] && f[185] && f[182];
	assign leaf[5622] = !f[332] && f[737] && !f[267];
	assign leaf[5623] = !f[332] && f[737] && f[267];
	assign leaf[5624] = f[332] && !f[371];
	assign leaf[5625] = f[332] && f[371];
	
	// Tree 385, Classifier 5, Iteration: 38
	assign leaf[5626] = !f[103] && !f[380] && !f[455] && !f[539];
	assign leaf[5627] = !f[103] && !f[380] && !f[455] && f[539];
	assign leaf[5628] = !f[103] && !f[380] && f[455] && !f[597];
	assign leaf[5629] = !f[103] && !f[380] && f[455] && f[597];
	assign leaf[5630] = !f[103] && f[380] && !f[325] && !f[243];
	assign leaf[5631] = !f[103] && f[380] && !f[325] && f[243];
	assign leaf[5632] = !f[103] && f[380] && f[325] && !f[321];
	assign leaf[5633] = !f[103] && f[380] && f[325] && f[321];
	assign leaf[5634] = f[103] && !f[243] && !f[324] && !f[319];
	assign leaf[5635] = f[103] && !f[243] && !f[324] && f[319];
	assign leaf[5636] = f[103] && !f[243] && f[324] && !f[437];
	assign leaf[5637] = f[103] && !f[243] && f[324] && f[437];
	assign leaf[5638] = f[103] && f[243];
	
	// Tree 386, Classifier 6, Iteration: 38
	assign leaf[5639] = !f[622] && !f[159] && !f[239] && !f[574];
	assign leaf[5640] = !f[622] && !f[159] && !f[239] && f[574];
	assign leaf[5641] = !f[622] && !f[159] && f[239] && !f[156];
	assign leaf[5642] = !f[622] && !f[159] && f[239] && f[156];
	assign leaf[5643] = !f[622] && f[159] && !f[325] && !f[328];
	assign leaf[5644] = !f[622] && f[159] && !f[325] && f[328];
	assign leaf[5645] = !f[622] && f[159] && f[325] && !f[467];
	assign leaf[5646] = !f[622] && f[159] && f[325] && f[467];
	assign leaf[5647] = f[622];
	
	// Tree 387, Classifier 7, Iteration: 38
	assign leaf[5648] = !f[122] && !f[160] && !f[129] && !f[325];
	assign leaf[5649] = !f[122] && !f[160] && !f[129] && f[325];
	assign leaf[5650] = !f[122] && !f[160] && f[129];
	assign leaf[5651] = !f[122] && f[160] && !f[684];
	assign leaf[5652] = !f[122] && f[160] && f[684];
	assign leaf[5653] = f[122];
	
	// Tree 388, Classifier 8, Iteration: 38
	assign leaf[5654] = !f[399] && !f[317] && !f[292] && !f[265];
	assign leaf[5655] = !f[399] && !f[317] && !f[292] && f[265];
	assign leaf[5656] = !f[399] && !f[317] && f[292] && !f[347];
	assign leaf[5657] = !f[399] && !f[317] && f[292] && f[347];
	assign leaf[5658] = !f[399] && f[317] && !f[290] && !f[372];
	assign leaf[5659] = !f[399] && f[317] && !f[290] && f[372];
	assign leaf[5660] = !f[399] && f[317] && f[290] && !f[517];
	assign leaf[5661] = !f[399] && f[317] && f[290] && f[517];
	assign leaf[5662] = f[399] && !f[607] && !f[304] && !f[287];
	assign leaf[5663] = f[399] && !f[607] && !f[304] && f[287];
	assign leaf[5664] = f[399] && !f[607] && f[304] && !f[212];
	assign leaf[5665] = f[399] && !f[607] && f[304] && f[212];
	assign leaf[5666] = f[399] && f[607] && !f[489] && !f[523];
	assign leaf[5667] = f[399] && f[607] && !f[489] && f[523];
	assign leaf[5668] = f[399] && f[607] && f[489] && !f[374];
	assign leaf[5669] = f[399] && f[607] && f[489] && f[374];
	
	// Tree 389, Classifier 9, Iteration: 38
	assign leaf[5670] = !f[368] && !f[437] && !f[549] && !f[382];
	assign leaf[5671] = !f[368] && !f[437] && !f[549] && f[382];
	assign leaf[5672] = !f[368] && !f[437] && f[549] && !f[462];
	assign leaf[5673] = !f[368] && !f[437] && f[549] && f[462];
	assign leaf[5674] = !f[368] && f[437] && !f[496] && !f[441];
	assign leaf[5675] = !f[368] && f[437] && !f[496] && f[441];
	assign leaf[5676] = !f[368] && f[437] && f[496] && !f[412];
	assign leaf[5677] = !f[368] && f[437] && f[496] && f[412];
	assign leaf[5678] = f[368] && !f[373] && !f[349] && !f[354];
	assign leaf[5679] = f[368] && !f[373] && !f[349] && f[354];
	assign leaf[5680] = f[368] && !f[373] && f[349];
	assign leaf[5681] = f[368] && f[373] && !f[465];
	assign leaf[5682] = f[368] && f[373] && f[465] && !f[260];
	assign leaf[5683] = f[368] && f[373] && f[465] && f[260];
	
	// Tree 390, Classifier 0, Iteration: 39
	assign leaf[5684] = !f[240] && !f[326] && !f[436] && !f[128];
	assign leaf[5685] = !f[240] && !f[326] && !f[436] && f[128];
	assign leaf[5686] = !f[240] && !f[326] && f[436] && !f[218];
	assign leaf[5687] = !f[240] && !f[326] && f[436] && f[218];
	assign leaf[5688] = !f[240] && f[326] && !f[236] && !f[381];
	assign leaf[5689] = !f[240] && f[326] && !f[236] && f[381];
	assign leaf[5690] = !f[240] && f[326] && f[236] && !f[397];
	assign leaf[5691] = !f[240] && f[326] && f[236] && f[397];
	assign leaf[5692] = f[240] && !f[326] && !f[538] && !f[466];
	assign leaf[5693] = f[240] && !f[326] && !f[538] && f[466];
	assign leaf[5694] = f[240] && !f[326] && f[538] && !f[608];
	assign leaf[5695] = f[240] && !f[326] && f[538] && f[608];
	assign leaf[5696] = f[240] && f[326] && !f[298] && !f[355];
	assign leaf[5697] = f[240] && f[326] && !f[298] && f[355];
	assign leaf[5698] = f[240] && f[326] && f[298] && !f[354];
	assign leaf[5699] = f[240] && f[326] && f[298] && f[354];
	
	// Tree 391, Classifier 1, Iteration: 39
	assign leaf[5700] = !f[683] && !f[95] && !f[314] && !f[609];
	assign leaf[5701] = !f[683] && !f[95] && !f[314] && f[609];
	assign leaf[5702] = !f[683] && !f[95] && f[314] && !f[184];
	assign leaf[5703] = !f[683] && !f[95] && f[314] && f[184];
	assign leaf[5704] = !f[683] && f[95] && !f[517];
	assign leaf[5705] = !f[683] && f[95] && f[517];
	assign leaf[5706] = f[683] && !f[268] && !f[185];
	assign leaf[5707] = f[683] && !f[268] && f[185];
	assign leaf[5708] = f[683] && f[268] && !f[208] && !f[347];
	assign leaf[5709] = f[683] && f[268] && !f[208] && f[347];
	assign leaf[5710] = f[683] && f[268] && f[208] && !f[319];
	assign leaf[5711] = f[683] && f[268] && f[208] && f[319];
	
	// Tree 392, Classifier 2, Iteration: 39
	assign leaf[5712] = !f[95] && !f[547] && !f[630] && !f[652];
	assign leaf[5713] = !f[95] && !f[547] && !f[630] && f[652];
	assign leaf[5714] = !f[95] && !f[547] && f[630] && !f[522];
	assign leaf[5715] = !f[95] && !f[547] && f[630] && f[522];
	assign leaf[5716] = !f[95] && f[547] && !f[685] && !f[687];
	assign leaf[5717] = !f[95] && f[547] && !f[685] && f[687];
	assign leaf[5718] = !f[95] && f[547] && f[685] && !f[461];
	assign leaf[5719] = !f[95] && f[547] && f[685] && f[461];
	assign leaf[5720] = f[95] && !f[354] && !f[458] && !f[461];
	assign leaf[5721] = f[95] && !f[354] && !f[458] && f[461];
	assign leaf[5722] = f[95] && !f[354] && f[458] && !f[517];
	assign leaf[5723] = f[95] && !f[354] && f[458] && f[517];
	assign leaf[5724] = f[95] && f[354] && !f[521];
	assign leaf[5725] = f[95] && f[354] && f[521] && !f[270];
	assign leaf[5726] = f[95] && f[354] && f[521] && f[270];
	
	// Tree 393, Classifier 3, Iteration: 39
	assign leaf[5727] = !f[358] && !f[486] && !f[456] && !f[595];
	assign leaf[5728] = !f[358] && !f[486] && !f[456] && f[595];
	assign leaf[5729] = !f[358] && !f[486] && f[456] && !f[299];
	assign leaf[5730] = !f[358] && !f[486] && f[456] && f[299];
	assign leaf[5731] = !f[358] && f[486] && !f[716] && !f[577];
	assign leaf[5732] = !f[358] && f[486] && !f[716] && f[577];
	assign leaf[5733] = !f[358] && f[486] && f[716] && !f[438];
	assign leaf[5734] = !f[358] && f[486] && f[716] && f[438];
	assign leaf[5735] = f[358] && !f[291] && !f[650];
	assign leaf[5736] = f[358] && !f[291] && f[650];
	assign leaf[5737] = f[358] && f[291] && !f[582] && !f[319];
	assign leaf[5738] = f[358] && f[291] && !f[582] && f[319];
	assign leaf[5739] = f[358] && f[291] && f[582];
	
	// Tree 394, Classifier 4, Iteration: 39
	assign leaf[5740] = !f[96] && !f[409] && !f[405] && !f[516];
	assign leaf[5741] = !f[96] && !f[409] && !f[405] && f[516];
	assign leaf[5742] = !f[96] && !f[409] && f[405] && !f[326];
	assign leaf[5743] = !f[96] && !f[409] && f[405] && f[326];
	assign leaf[5744] = !f[96] && f[409] && !f[375] && !f[293];
	assign leaf[5745] = !f[96] && f[409] && !f[375] && f[293];
	assign leaf[5746] = !f[96] && f[409] && f[375] && !f[241];
	assign leaf[5747] = !f[96] && f[409] && f[375] && f[241];
	assign leaf[5748] = f[96] && !f[574];
	assign leaf[5749] = f[96] && f[574];
	
	// Tree 395, Classifier 5, Iteration: 39
	assign leaf[5750] = !f[304] && !f[188] && !f[490] && !f[239];
	assign leaf[5751] = !f[304] && !f[188] && !f[490] && f[239];
	assign leaf[5752] = !f[304] && !f[188] && f[490] && !f[273];
	assign leaf[5753] = !f[304] && !f[188] && f[490] && f[273];
	assign leaf[5754] = !f[304] && f[188] && !f[212] && !f[216];
	assign leaf[5755] = !f[304] && f[188] && !f[212] && f[216];
	assign leaf[5756] = !f[304] && f[188] && f[212] && !f[300];
	assign leaf[5757] = !f[304] && f[188] && f[212] && f[300];
	assign leaf[5758] = f[304] && !f[301] && !f[217];
	assign leaf[5759] = f[304] && !f[301] && f[217];
	assign leaf[5760] = f[304] && f[301] && !f[383] && !f[234];
	assign leaf[5761] = f[304] && f[301] && !f[383] && f[234];
	assign leaf[5762] = f[304] && f[301] && f[383];
	
	// Tree 396, Classifier 6, Iteration: 39
	assign leaf[5763] = !f[91] && !f[682] && !f[459] && !f[457];
	assign leaf[5764] = !f[91] && !f[682] && !f[459] && f[457];
	assign leaf[5765] = !f[91] && !f[682] && f[459] && !f[403];
	assign leaf[5766] = !f[91] && !f[682] && f[459] && f[403];
	assign leaf[5767] = !f[91] && f[682];
	assign leaf[5768] = f[91] && !f[356];
	assign leaf[5769] = f[91] && f[356];
	
	// Tree 397, Classifier 7, Iteration: 39
	assign leaf[5770] = !f[124] && !f[459] && !f[183] && !f[151];
	assign leaf[5771] = !f[124] && !f[459] && !f[183] && f[151];
	assign leaf[5772] = !f[124] && !f[459] && f[183] && !f[321];
	assign leaf[5773] = !f[124] && !f[459] && f[183] && f[321];
	assign leaf[5774] = !f[124] && f[459] && !f[400] && !f[324];
	assign leaf[5775] = !f[124] && f[459] && !f[400] && f[324];
	assign leaf[5776] = !f[124] && f[459] && f[400] && !f[469];
	assign leaf[5777] = !f[124] && f[459] && f[400] && f[469];
	assign leaf[5778] = f[124];
	
	// Tree 398, Classifier 8, Iteration: 39
	assign leaf[5779] = !f[219] && !f[412] && !f[688] && !f[350];
	assign leaf[5780] = !f[219] && !f[412] && !f[688] && f[350];
	assign leaf[5781] = !f[219] && !f[412] && f[688] && !f[545];
	assign leaf[5782] = !f[219] && !f[412] && f[688] && f[545];
	assign leaf[5783] = !f[219] && f[412] && !f[332] && !f[126];
	assign leaf[5784] = !f[219] && f[412] && !f[332] && f[126];
	assign leaf[5785] = !f[219] && f[412] && f[332] && !f[344];
	assign leaf[5786] = !f[219] && f[412] && f[332] && f[344];
	assign leaf[5787] = f[219] && !f[454] && !f[649] && !f[379];
	assign leaf[5788] = f[219] && !f[454] && !f[649] && f[379];
	assign leaf[5789] = f[219] && !f[454] && f[649] && !f[597];
	assign leaf[5790] = f[219] && !f[454] && f[649] && f[597];
	assign leaf[5791] = f[219] && f[454] && !f[272] && !f[181];
	assign leaf[5792] = f[219] && f[454] && !f[272] && f[181];
	assign leaf[5793] = f[219] && f[454] && f[272] && !f[595];
	assign leaf[5794] = f[219] && f[454] && f[272] && f[595];
	
	// Tree 399, Classifier 9, Iteration: 39
	assign leaf[5795] = !f[350] && !f[486] && !f[406] && !f[512];
	assign leaf[5796] = !f[350] && !f[486] && !f[406] && f[512];
	assign leaf[5797] = !f[350] && !f[486] && f[406] && !f[489];
	assign leaf[5798] = !f[350] && !f[486] && f[406] && f[489];
	assign leaf[5799] = !f[350] && f[486] && !f[431] && !f[428];
	assign leaf[5800] = !f[350] && f[486] && !f[431] && f[428];
	assign leaf[5801] = !f[350] && f[486] && f[431] && !f[428];
	assign leaf[5802] = !f[350] && f[486] && f[431] && f[428];
	assign leaf[5803] = f[350] && !f[325] && !f[434] && !f[464];
	assign leaf[5804] = f[350] && !f[325] && !f[434] && f[464];
	assign leaf[5805] = f[350] && !f[325] && f[434] && !f[264];
	assign leaf[5806] = f[350] && !f[325] && f[434] && f[264];
	assign leaf[5807] = f[350] && f[325] && !f[460] && !f[456];
	assign leaf[5808] = f[350] && f[325] && !f[460] && f[456];
	assign leaf[5809] = f[350] && f[325] && f[460] && !f[345];
	assign leaf[5810] = f[350] && f[325] && f[460] && f[345];
	
	// Tree 400, Classifier 0, Iteration: 40
	assign leaf[5811] = !f[688] && !f[453] && !f[298] && !f[300];
	assign leaf[5812] = !f[688] && !f[453] && !f[298] && f[300];
	assign leaf[5813] = !f[688] && !f[453] && f[298] && !f[459];
	assign leaf[5814] = !f[688] && !f[453] && f[298] && f[459];
	assign leaf[5815] = !f[688] && f[453] && !f[459] && !f[383];
	assign leaf[5816] = !f[688] && f[453] && !f[459] && f[383];
	assign leaf[5817] = !f[688] && f[453] && f[459] && !f[572];
	assign leaf[5818] = !f[688] && f[453] && f[459] && f[572];
	assign leaf[5819] = f[688] && !f[657] && !f[549];
	assign leaf[5820] = f[688] && !f[657] && f[549] && !f[273];
	assign leaf[5821] = f[688] && !f[657] && f[549] && f[273];
	assign leaf[5822] = f[688] && f[657] && !f[186] && !f[655];
	assign leaf[5823] = f[688] && f[657] && !f[186] && f[655];
	assign leaf[5824] = f[688] && f[657] && f[186] && !f[272];
	assign leaf[5825] = f[688] && f[657] && f[186] && f[272];
	
	// Tree 401, Classifier 1, Iteration: 40
	assign leaf[5826] = !f[468] && !f[716] && !f[680] && !f[685];
	assign leaf[5827] = !f[468] && !f[716] && !f[680] && f[685];
	assign leaf[5828] = !f[468] && !f[716] && f[680] && !f[211];
	assign leaf[5829] = !f[468] && !f[716] && f[680] && f[211];
	assign leaf[5830] = !f[468] && f[716];
	assign leaf[5831] = f[468];
	
	// Tree 402, Classifier 2, Iteration: 40
	assign leaf[5832] = !f[666] && !f[611] && !f[556] && !f[472];
	assign leaf[5833] = !f[666] && !f[611] && !f[556] && f[472];
	assign leaf[5834] = !f[666] && !f[611] && f[556] && !f[127];
	assign leaf[5835] = !f[666] && !f[611] && f[556] && f[127];
	assign leaf[5836] = !f[666] && f[611] && !f[527] && !f[344];
	assign leaf[5837] = !f[666] && f[611] && !f[527] && f[344];
	assign leaf[5838] = !f[666] && f[611] && f[527] && !f[293];
	assign leaf[5839] = !f[666] && f[611] && f[527] && f[293];
	assign leaf[5840] = f[666] && !f[525] && !f[582] && !f[576];
	assign leaf[5841] = f[666] && !f[525] && !f[582] && f[576];
	assign leaf[5842] = f[666] && !f[525] && f[582];
	assign leaf[5843] = f[666] && f[525] && !f[155];
	assign leaf[5844] = f[666] && f[525] && f[155];
	
	// Tree 403, Classifier 3, Iteration: 40
	assign leaf[5845] = !f[210] && !f[234] && !f[156] && !f[525];
	assign leaf[5846] = !f[210] && !f[234] && !f[156] && f[525];
	assign leaf[5847] = !f[210] && !f[234] && f[156] && !f[236];
	assign leaf[5848] = !f[210] && !f[234] && f[156] && f[236];
	assign leaf[5849] = !f[210] && f[234] && !f[151] && !f[491];
	assign leaf[5850] = !f[210] && f[234] && !f[151] && f[491];
	assign leaf[5851] = !f[210] && f[234] && f[151] && !f[258];
	assign leaf[5852] = !f[210] && f[234] && f[151] && f[258];
	assign leaf[5853] = f[210] && !f[346] && !f[572] && !f[489];
	assign leaf[5854] = f[210] && !f[346] && !f[572] && f[489];
	assign leaf[5855] = f[210] && !f[346] && f[572] && !f[536];
	assign leaf[5856] = f[210] && !f[346] && f[572] && f[536];
	assign leaf[5857] = f[210] && f[346] && !f[442] && !f[375];
	assign leaf[5858] = f[210] && f[346] && !f[442] && f[375];
	assign leaf[5859] = f[210] && f[346] && f[442] && !f[314];
	assign leaf[5860] = f[210] && f[346] && f[442] && f[314];
	
	// Tree 404, Classifier 4, Iteration: 40
	assign leaf[5861] = !f[465] && !f[605] && !f[238] && !f[294];
	assign leaf[5862] = !f[465] && !f[605] && !f[238] && f[294];
	assign leaf[5863] = !f[465] && !f[605] && f[238] && !f[240];
	assign leaf[5864] = !f[465] && !f[605] && f[238] && f[240];
	assign leaf[5865] = !f[465] && f[605] && !f[218] && !f[662];
	assign leaf[5866] = !f[465] && f[605] && !f[218] && f[662];
	assign leaf[5867] = !f[465] && f[605] && f[218] && !f[291];
	assign leaf[5868] = !f[465] && f[605] && f[218] && f[291];
	assign leaf[5869] = f[465] && !f[381] && !f[297] && !f[214];
	assign leaf[5870] = f[465] && !f[381] && !f[297] && f[214];
	assign leaf[5871] = f[465] && !f[381] && f[297] && !f[549];
	assign leaf[5872] = f[465] && !f[381] && f[297] && f[549];
	assign leaf[5873] = f[465] && f[381] && !f[375] && !f[355];
	assign leaf[5874] = f[465] && f[381] && !f[375] && f[355];
	assign leaf[5875] = f[465] && f[381] && f[375] && !f[715];
	assign leaf[5876] = f[465] && f[381] && f[375] && f[715];
	
	// Tree 405, Classifier 5, Iteration: 40
	assign leaf[5877] = !f[276] && !f[200] && !f[332] && !f[329];
	assign leaf[5878] = !f[276] && !f[200] && !f[332] && f[329];
	assign leaf[5879] = !f[276] && !f[200] && f[332] && !f[214];
	assign leaf[5880] = !f[276] && !f[200] && f[332] && f[214];
	assign leaf[5881] = !f[276] && f[200] && !f[236];
	assign leaf[5882] = !f[276] && f[200] && f[236];
	assign leaf[5883] = f[276] && !f[186] && !f[357] && !f[180];
	assign leaf[5884] = f[276] && !f[186] && !f[357] && f[180];
	assign leaf[5885] = f[276] && !f[186] && f[357];
	assign leaf[5886] = f[276] && f[186] && !f[244];
	assign leaf[5887] = f[276] && f[186] && f[244];
	
	// Tree 406, Classifier 6, Iteration: 40
	assign leaf[5888] = !f[609] && !f[93] && !f[270] && !f[274];
	assign leaf[5889] = !f[609] && !f[93] && !f[270] && f[274];
	assign leaf[5890] = !f[609] && !f[93] && f[270] && !f[350];
	assign leaf[5891] = !f[609] && !f[93] && f[270] && f[350];
	assign leaf[5892] = !f[609] && f[93] && !f[123] && !f[431];
	assign leaf[5893] = !f[609] && f[93] && !f[123] && f[431];
	assign leaf[5894] = !f[609] && f[93] && f[123] && !f[206];
	assign leaf[5895] = !f[609] && f[93] && f[123] && f[206];
	assign leaf[5896] = f[609] && !f[455] && !f[551] && !f[290];
	assign leaf[5897] = f[609] && !f[455] && !f[551] && f[290];
	assign leaf[5898] = f[609] && !f[455] && f[551] && !f[555];
	assign leaf[5899] = f[609] && !f[455] && f[551] && f[555];
	assign leaf[5900] = f[609] && f[455] && !f[633] && !f[573];
	assign leaf[5901] = f[609] && f[455] && !f[633] && f[573];
	assign leaf[5902] = f[609] && f[455] && f[633] && !f[205];
	assign leaf[5903] = f[609] && f[455] && f[633] && f[205];
	
	// Tree 407, Classifier 7, Iteration: 40
	assign leaf[5904] = !f[510] && !f[411] && !f[242] && !f[467];
	assign leaf[5905] = !f[510] && !f[411] && !f[242] && f[467];
	assign leaf[5906] = !f[510] && !f[411] && f[242] && !f[578];
	assign leaf[5907] = !f[510] && !f[411] && f[242] && f[578];
	assign leaf[5908] = !f[510] && f[411] && !f[383] && !f[551];
	assign leaf[5909] = !f[510] && f[411] && !f[383] && f[551];
	assign leaf[5910] = !f[510] && f[411] && f[383] && !f[460];
	assign leaf[5911] = !f[510] && f[411] && f[383] && f[460];
	assign leaf[5912] = f[510] && !f[257] && !f[541] && !f[519];
	assign leaf[5913] = f[510] && !f[257] && !f[541] && f[519];
	assign leaf[5914] = f[510] && !f[257] && f[541] && !f[219];
	assign leaf[5915] = f[510] && !f[257] && f[541] && f[219];
	assign leaf[5916] = f[510] && f[257];
	
	// Tree 408, Classifier 8, Iteration: 40
	assign leaf[5917] = !f[340] && !f[468] && !f[357] && !f[410];
	assign leaf[5918] = !f[340] && !f[468] && !f[357] && f[410];
	assign leaf[5919] = !f[340] && !f[468] && f[357] && !f[326];
	assign leaf[5920] = !f[340] && !f[468] && f[357] && f[326];
	assign leaf[5921] = !f[340] && f[468] && !f[577] && !f[492];
	assign leaf[5922] = !f[340] && f[468] && !f[577] && f[492];
	assign leaf[5923] = !f[340] && f[468] && f[577] && !f[380];
	assign leaf[5924] = !f[340] && f[468] && f[577] && f[380];
	assign leaf[5925] = f[340] && !f[464];
	assign leaf[5926] = f[340] && f[464] && !f[152] && !f[321];
	assign leaf[5927] = f[340] && f[464] && !f[152] && f[321];
	assign leaf[5928] = f[340] && f[464] && f[152];
	
	// Tree 409, Classifier 9, Iteration: 40
	assign leaf[5929] = !f[408] && !f[439] && !f[410] && !f[550];
	assign leaf[5930] = !f[408] && !f[439] && !f[410] && f[550];
	assign leaf[5931] = !f[408] && !f[439] && f[410] && !f[324];
	assign leaf[5932] = !f[408] && !f[439] && f[410] && f[324];
	assign leaf[5933] = !f[408] && f[439] && !f[373] && !f[207];
	assign leaf[5934] = !f[408] && f[439] && !f[373] && f[207];
	assign leaf[5935] = !f[408] && f[439] && f[373] && !f[155];
	assign leaf[5936] = !f[408] && f[439] && f[373] && f[155];
	assign leaf[5937] = f[408] && !f[149] && !f[517] && !f[181];
	assign leaf[5938] = f[408] && !f[149] && !f[517] && f[181];
	assign leaf[5939] = f[408] && !f[149] && f[517] && !f[630];
	assign leaf[5940] = f[408] && !f[149] && f[517] && f[630];
	assign leaf[5941] = f[408] && f[149] && !f[286];
	assign leaf[5942] = f[408] && f[149] && f[286];
	
	// Tree 410, Classifier 0, Iteration: 41
	assign leaf[5943] = !f[444] && !f[319] && !f[494] && !f[413];
	assign leaf[5944] = !f[444] && !f[319] && !f[494] && f[413];
	assign leaf[5945] = !f[444] && !f[319] && f[494] && !f[657];
	assign leaf[5946] = !f[444] && !f[319] && f[494] && f[657];
	assign leaf[5947] = !f[444] && f[319] && !f[605] && !f[493];
	assign leaf[5948] = !f[444] && f[319] && !f[605] && f[493];
	assign leaf[5949] = !f[444] && f[319] && f[605] && !f[320];
	assign leaf[5950] = !f[444] && f[319] && f[605] && f[320];
	assign leaf[5951] = f[444] && !f[152] && !f[289];
	assign leaf[5952] = f[444] && !f[152] && f[289] && !f[600];
	assign leaf[5953] = f[444] && !f[152] && f[289] && f[600];
	assign leaf[5954] = f[444] && f[152] && !f[483];
	assign leaf[5955] = f[444] && f[152] && f[483] && !f[302];
	assign leaf[5956] = f[444] && f[152] && f[483] && f[302];
	
	// Tree 411, Classifier 1, Iteration: 41
	assign leaf[5957] = !f[383] && !f[518] && !f[631] && !f[210];
	assign leaf[5958] = !f[383] && !f[518] && !f[631] && f[210];
	assign leaf[5959] = !f[383] && !f[518] && f[631] && !f[405];
	assign leaf[5960] = !f[383] && !f[518] && f[631] && f[405];
	assign leaf[5961] = !f[383] && f[518] && !f[603] && !f[181];
	assign leaf[5962] = !f[383] && f[518] && !f[603] && f[181];
	assign leaf[5963] = !f[383] && f[518] && f[603] && !f[573];
	assign leaf[5964] = !f[383] && f[518] && f[603] && f[573];
	assign leaf[5965] = f[383] && !f[300] && !f[380];
	assign leaf[5966] = f[383] && !f[300] && f[380];
	assign leaf[5967] = f[383] && f[300] && !f[213];
	assign leaf[5968] = f[383] && f[300] && f[213];
	
	// Tree 412, Classifier 2, Iteration: 41
	assign leaf[5969] = !f[409] && !f[354] && !f[97] && !f[149];
	assign leaf[5970] = !f[409] && !f[354] && !f[97] && f[149];
	assign leaf[5971] = !f[409] && !f[354] && f[97] && !f[463];
	assign leaf[5972] = !f[409] && !f[354] && f[97] && f[463];
	assign leaf[5973] = !f[409] && f[354] && !f[294] && !f[210];
	assign leaf[5974] = !f[409] && f[354] && !f[294] && f[210];
	assign leaf[5975] = !f[409] && f[354] && f[294] && !f[371];
	assign leaf[5976] = !f[409] && f[354] && f[294] && f[371];
	assign leaf[5977] = f[409] && !f[463] && !f[355] && !f[379];
	assign leaf[5978] = f[409] && !f[463] && !f[355] && f[379];
	assign leaf[5979] = f[409] && !f[463] && f[355] && !f[655];
	assign leaf[5980] = f[409] && !f[463] && f[355] && f[655];
	assign leaf[5981] = f[409] && f[463] && !f[538] && !f[460];
	assign leaf[5982] = f[409] && f[463] && !f[538] && f[460];
	assign leaf[5983] = f[409] && f[463] && f[538] && !f[600];
	assign leaf[5984] = f[409] && f[463] && f[538] && f[600];
	
	// Tree 413, Classifier 3, Iteration: 41
	assign leaf[5985] = !f[269] && !f[513] && !f[497] && !f[299];
	assign leaf[5986] = !f[269] && !f[513] && !f[497] && f[299];
	assign leaf[5987] = !f[269] && !f[513] && f[497] && !f[265];
	assign leaf[5988] = !f[269] && !f[513] && f[497] && f[265];
	assign leaf[5989] = !f[269] && f[513] && !f[509] && !f[523];
	assign leaf[5990] = !f[269] && f[513] && !f[509] && f[523];
	assign leaf[5991] = !f[269] && f[513] && f[509] && !f[462];
	assign leaf[5992] = !f[269] && f[513] && f[509] && f[462];
	assign leaf[5993] = f[269] && !f[341] && !f[323] && !f[433];
	assign leaf[5994] = f[269] && !f[341] && !f[323] && f[433];
	assign leaf[5995] = f[269] && !f[341] && f[323] && !f[494];
	assign leaf[5996] = f[269] && !f[341] && f[323] && f[494];
	assign leaf[5997] = f[269] && f[341] && !f[656];
	assign leaf[5998] = f[269] && f[341] && f[656] && !f[399];
	assign leaf[5999] = f[269] && f[341] && f[656] && f[399];
	
	// Tree 414, Classifier 4, Iteration: 41
	assign leaf[6000] = !f[96] && !f[346] && !f[625] && !f[348];
	assign leaf[6001] = !f[96] && !f[346] && !f[625] && f[348];
	assign leaf[6002] = !f[96] && !f[346] && f[625] && !f[709];
	assign leaf[6003] = !f[96] && !f[346] && f[625] && f[709];
	assign leaf[6004] = !f[96] && f[346] && !f[340] && !f[400];
	assign leaf[6005] = !f[96] && f[346] && !f[340] && f[400];
	assign leaf[6006] = !f[96] && f[346] && f[340] && !f[398];
	assign leaf[6007] = !f[96] && f[346] && f[340] && f[398];
	assign leaf[6008] = f[96] && !f[455];
	assign leaf[6009] = f[96] && f[455];
	
	// Tree 415, Classifier 5, Iteration: 41
	assign leaf[6010] = !f[103] && !f[436] && !f[485] && !f[402];
	assign leaf[6011] = !f[103] && !f[436] && !f[485] && f[402];
	assign leaf[6012] = !f[103] && !f[436] && f[485] && !f[541];
	assign leaf[6013] = !f[103] && !f[436] && f[485] && f[541];
	assign leaf[6014] = !f[103] && f[436] && !f[354] && !f[215];
	assign leaf[6015] = !f[103] && f[436] && !f[354] && f[215];
	assign leaf[6016] = !f[103] && f[436] && f[354] && !f[321];
	assign leaf[6017] = !f[103] && f[436] && f[354] && f[321];
	assign leaf[6018] = f[103] && !f[245] && !f[576];
	assign leaf[6019] = f[103] && !f[245] && f[576] && !f[348];
	assign leaf[6020] = f[103] && !f[245] && f[576] && f[348];
	assign leaf[6021] = f[103] && f[245];
	
	// Tree 416, Classifier 6, Iteration: 41
	assign leaf[6022] = !f[622] && !f[208] && !f[98] && !f[550];
	assign leaf[6023] = !f[622] && !f[208] && !f[98] && f[550];
	assign leaf[6024] = !f[622] && !f[208] && f[98] && !f[551];
	assign leaf[6025] = !f[622] && !f[208] && f[98] && f[551];
	assign leaf[6026] = !f[622] && f[208] && !f[318] && !f[416];
	assign leaf[6027] = !f[622] && f[208] && !f[318] && f[416];
	assign leaf[6028] = !f[622] && f[208] && f[318] && !f[178];
	assign leaf[6029] = !f[622] && f[208] && f[318] && f[178];
	assign leaf[6030] = f[622];
	
	// Tree 417, Classifier 7, Iteration: 41
	assign leaf[6031] = !f[158] && !f[637] && !f[202] && !f[549];
	assign leaf[6032] = !f[158] && !f[637] && !f[202] && f[549];
	assign leaf[6033] = !f[158] && !f[637] && f[202] && !f[493];
	assign leaf[6034] = !f[158] && !f[637] && f[202] && f[493];
	assign leaf[6035] = !f[158] && f[637] && !f[318];
	assign leaf[6036] = !f[158] && f[637] && f[318] && !f[179];
	assign leaf[6037] = !f[158] && f[637] && f[318] && f[179];
	assign leaf[6038] = f[158] && !f[154] && !f[232] && !f[377];
	assign leaf[6039] = f[158] && !f[154] && !f[232] && f[377];
	assign leaf[6040] = f[158] && !f[154] && f[232];
	assign leaf[6041] = f[158] && f[154] && !f[235];
	assign leaf[6042] = f[158] && f[154] && f[235] && !f[263];
	assign leaf[6043] = f[158] && f[154] && f[235] && f[263];
	
	// Tree 418, Classifier 8, Iteration: 41
	assign leaf[6044] = !f[437] && !f[492] && !f[547] && !f[543];
	assign leaf[6045] = !f[437] && !f[492] && !f[547] && f[543];
	assign leaf[6046] = !f[437] && !f[492] && f[547] && !f[550];
	assign leaf[6047] = !f[437] && !f[492] && f[547] && f[550];
	assign leaf[6048] = !f[437] && f[492] && !f[406] && !f[219];
	assign leaf[6049] = !f[437] && f[492] && !f[406] && f[219];
	assign leaf[6050] = !f[437] && f[492] && f[406] && !f[518];
	assign leaf[6051] = !f[437] && f[492] && f[406] && f[518];
	assign leaf[6052] = f[437] && !f[353] && !f[489] && !f[323];
	assign leaf[6053] = f[437] && !f[353] && !f[489] && f[323];
	assign leaf[6054] = f[437] && !f[353] && f[489] && !f[483];
	assign leaf[6055] = f[437] && !f[353] && f[489] && f[483];
	assign leaf[6056] = f[437] && f[353] && !f[491] && !f[483];
	assign leaf[6057] = f[437] && f[353] && !f[491] && f[483];
	assign leaf[6058] = f[437] && f[353] && f[491] && !f[662];
	assign leaf[6059] = f[437] && f[353] && f[491] && f[662];
	
	// Tree 419, Classifier 9, Iteration: 41
	assign leaf[6060] = !f[500] && !f[273] && !f[327] && !f[439];
	assign leaf[6061] = !f[500] && !f[273] && !f[327] && f[439];
	assign leaf[6062] = !f[500] && !f[273] && f[327] && !f[351];
	assign leaf[6063] = !f[500] && !f[273] && f[327] && f[351];
	assign leaf[6064] = !f[500] && f[273] && !f[215] && !f[241];
	assign leaf[6065] = !f[500] && f[273] && !f[215] && f[241];
	assign leaf[6066] = !f[500] && f[273] && f[215] && !f[385];
	assign leaf[6067] = !f[500] && f[273] && f[215] && f[385];
	assign leaf[6068] = f[500] && !f[416];
	assign leaf[6069] = f[500] && f[416];
	
	// Tree 420, Classifier 0, Iteration: 42
	assign leaf[6070] = !f[347] && !f[466] && !f[404] && !f[293];
	assign leaf[6071] = !f[347] && !f[466] && !f[404] && f[293];
	assign leaf[6072] = !f[347] && !f[466] && f[404] && !f[465];
	assign leaf[6073] = !f[347] && !f[466] && f[404] && f[465];
	assign leaf[6074] = !f[347] && f[466] && !f[127] && !f[329];
	assign leaf[6075] = !f[347] && f[466] && !f[127] && f[329];
	assign leaf[6076] = !f[347] && f[466] && f[127] && !f[344];
	assign leaf[6077] = !f[347] && f[466] && f[127] && f[344];
	assign leaf[6078] = f[347] && !f[493] && !f[348] && !f[551];
	assign leaf[6079] = f[347] && !f[493] && !f[348] && f[551];
	assign leaf[6080] = f[347] && !f[493] && f[348] && !f[273];
	assign leaf[6081] = f[347] && !f[493] && f[348] && f[273];
	assign leaf[6082] = f[347] && f[493] && !f[577] && !f[523];
	assign leaf[6083] = f[347] && f[493] && !f[577] && f[523];
	assign leaf[6084] = f[347] && f[493] && f[577] && !f[491];
	assign leaf[6085] = f[347] && f[493] && f[577] && f[491];
	
	// Tree 421, Classifier 1, Iteration: 42
	assign leaf[6086] = !f[244] && !f[293] && !f[181] && !f[604];
	assign leaf[6087] = !f[244] && !f[293] && !f[181] && f[604];
	assign leaf[6088] = !f[244] && !f[293] && f[181] && !f[405];
	assign leaf[6089] = !f[244] && !f[293] && f[181] && f[405];
	assign leaf[6090] = !f[244] && f[293] && !f[160] && !f[321];
	assign leaf[6091] = !f[244] && f[293] && !f[160] && f[321];
	assign leaf[6092] = !f[244] && f[293] && f[160] && !f[238];
	assign leaf[6093] = !f[244] && f[293] && f[160] && f[238];
	assign leaf[6094] = f[244] && !f[265] && !f[156] && !f[325];
	assign leaf[6095] = f[244] && !f[265] && !f[156] && f[325];
	assign leaf[6096] = f[244] && !f[265] && f[156] && !f[404];
	assign leaf[6097] = f[244] && !f[265] && f[156] && f[404];
	assign leaf[6098] = f[244] && f[265] && !f[577] && !f[291];
	assign leaf[6099] = f[244] && f[265] && !f[577] && f[291];
	assign leaf[6100] = f[244] && f[265] && f[577];
	
	// Tree 422, Classifier 2, Iteration: 42
	assign leaf[6101] = !f[409] && !f[549] && !f[605] && !f[443];
	assign leaf[6102] = !f[409] && !f[549] && !f[605] && f[443];
	assign leaf[6103] = !f[409] && !f[549] && f[605] && !f[523];
	assign leaf[6104] = !f[409] && !f[549] && f[605] && f[523];
	assign leaf[6105] = !f[409] && f[549] && !f[660] && !f[460];
	assign leaf[6106] = !f[409] && f[549] && !f[660] && f[460];
	assign leaf[6107] = !f[409] && f[549] && f[660] && !f[384];
	assign leaf[6108] = !f[409] && f[549] && f[660] && f[384];
	assign leaf[6109] = f[409] && !f[463] && !f[176] && !f[681];
	assign leaf[6110] = f[409] && !f[463] && !f[176] && f[681];
	assign leaf[6111] = f[409] && !f[463] && f[176] && !f[521];
	assign leaf[6112] = f[409] && !f[463] && f[176] && f[521];
	assign leaf[6113] = f[409] && f[463] && !f[609] && !f[201];
	assign leaf[6114] = f[409] && f[463] && !f[609] && f[201];
	assign leaf[6115] = f[409] && f[463] && f[609] && !f[469];
	assign leaf[6116] = f[409] && f[463] && f[609] && f[469];
	
	// Tree 423, Classifier 3, Iteration: 42
	assign leaf[6117] = !f[371] && !f[211] && !f[235] && !f[156];
	assign leaf[6118] = !f[371] && !f[211] && !f[235] && f[156];
	assign leaf[6119] = !f[371] && !f[211] && f[235] && !f[202];
	assign leaf[6120] = !f[371] && !f[211] && f[235] && f[202];
	assign leaf[6121] = !f[371] && f[211] && !f[131] && !f[549];
	assign leaf[6122] = !f[371] && f[211] && !f[131] && f[549];
	assign leaf[6123] = !f[371] && f[211] && f[131] && !f[266];
	assign leaf[6124] = !f[371] && f[211] && f[131] && f[266];
	assign leaf[6125] = f[371] && !f[315] && !f[313] && !f[481];
	assign leaf[6126] = f[371] && !f[315] && !f[313] && f[481];
	assign leaf[6127] = f[371] && !f[315] && f[313];
	assign leaf[6128] = f[371] && f[315] && !f[232] && !f[351];
	assign leaf[6129] = f[371] && f[315] && !f[232] && f[351];
	assign leaf[6130] = f[371] && f[315] && f[232] && !f[689];
	assign leaf[6131] = f[371] && f[315] && f[232] && f[689];
	
	// Tree 424, Classifier 4, Iteration: 42
	assign leaf[6132] = !f[625] && !f[491] && !f[321] && !f[411];
	assign leaf[6133] = !f[625] && !f[491] && !f[321] && f[411];
	assign leaf[6134] = !f[625] && !f[491] && f[321] && !f[654];
	assign leaf[6135] = !f[625] && !f[491] && f[321] && f[654];
	assign leaf[6136] = !f[625] && f[491] && !f[326] && !f[243];
	assign leaf[6137] = !f[625] && f[491] && !f[326] && f[243];
	assign leaf[6138] = !f[625] && f[491] && f[326] && !f[379];
	assign leaf[6139] = !f[625] && f[491] && f[326] && f[379];
	assign leaf[6140] = f[625] && !f[543] && !f[190];
	assign leaf[6141] = f[625] && !f[543] && f[190] && !f[596];
	assign leaf[6142] = f[625] && !f[543] && f[190] && f[596];
	assign leaf[6143] = f[625] && f[543] && !f[186] && !f[268];
	assign leaf[6144] = f[625] && f[543] && !f[186] && f[268];
	assign leaf[6145] = f[625] && f[543] && f[186] && !f[132];
	assign leaf[6146] = f[625] && f[543] && f[186] && f[132];
	
	// Tree 425, Classifier 5, Iteration: 42
	assign leaf[6147] = !f[612] && !f[565] && !f[289] && !f[481];
	assign leaf[6148] = !f[612] && !f[565] && !f[289] && f[481];
	assign leaf[6149] = !f[612] && !f[565] && f[289] && !f[205];
	assign leaf[6150] = !f[612] && !f[565] && f[289] && f[205];
	assign leaf[6151] = !f[612] && f[565] && !f[454] && !f[294];
	assign leaf[6152] = !f[612] && f[565] && !f[454] && f[294];
	assign leaf[6153] = !f[612] && f[565] && f[454] && !f[246];
	assign leaf[6154] = !f[612] && f[565] && f[454] && f[246];
	assign leaf[6155] = f[612];
	
	// Tree 426, Classifier 6, Iteration: 42
	assign leaf[6156] = !f[594] && !f[685] && !f[661] && !f[635];
	assign leaf[6157] = !f[594] && !f[685] && !f[661] && f[635];
	assign leaf[6158] = !f[594] && !f[685] && f[661] && !f[158];
	assign leaf[6159] = !f[594] && !f[685] && f[661] && f[158];
	assign leaf[6160] = !f[594] && f[685] && !f[598];
	assign leaf[6161] = !f[594] && f[685] && f[598] && !f[381];
	assign leaf[6162] = !f[594] && f[685] && f[598] && f[381];
	assign leaf[6163] = f[594] && !f[400] && !f[185] && !f[543];
	assign leaf[6164] = f[594] && !f[400] && !f[185] && f[543];
	assign leaf[6165] = f[594] && !f[400] && f[185];
	assign leaf[6166] = f[594] && f[400] && !f[217] && !f[435];
	assign leaf[6167] = f[594] && f[400] && !f[217] && f[435];
	assign leaf[6168] = f[594] && f[400] && f[217];
	
	// Tree 427, Classifier 7, Iteration: 42
	assign leaf[6169] = !f[677] && !f[595] && !f[434] && !f[378];
	assign leaf[6170] = !f[677] && !f[595] && !f[434] && f[378];
	assign leaf[6171] = !f[677] && !f[595] && f[434] && !f[351];
	assign leaf[6172] = !f[677] && !f[595] && f[434] && f[351];
	assign leaf[6173] = !f[677] && f[595] && !f[573] && !f[656];
	assign leaf[6174] = !f[677] && f[595] && !f[573] && f[656];
	assign leaf[6175] = !f[677] && f[595] && f[573];
	assign leaf[6176] = f[677] && !f[404] && !f[681] && !f[234];
	assign leaf[6177] = f[677] && !f[404] && !f[681] && f[234];
	assign leaf[6178] = f[677] && !f[404] && f[681];
	assign leaf[6179] = f[677] && f[404];
	
	// Tree 428, Classifier 8, Iteration: 42
	assign leaf[6180] = !f[303] && !f[650] && !f[244] && !f[637];
	assign leaf[6181] = !f[303] && !f[650] && !f[244] && f[637];
	assign leaf[6182] = !f[303] && !f[650] && f[244] && !f[242];
	assign leaf[6183] = !f[303] && !f[650] && f[244] && f[242];
	assign leaf[6184] = !f[303] && f[650] && !f[539] && !f[541];
	assign leaf[6185] = !f[303] && f[650] && !f[539] && f[541];
	assign leaf[6186] = !f[303] && f[650] && f[539] && !f[634];
	assign leaf[6187] = !f[303] && f[650] && f[539] && f[634];
	assign leaf[6188] = f[303] && !f[485] && !f[577] && !f[301];
	assign leaf[6189] = f[303] && !f[485] && !f[577] && f[301];
	assign leaf[6190] = f[303] && !f[485] && f[577] && !f[409];
	assign leaf[6191] = f[303] && !f[485] && f[577] && f[409];
	assign leaf[6192] = f[303] && f[485] && !f[207] && !f[492];
	assign leaf[6193] = f[303] && f[485] && !f[207] && f[492];
	assign leaf[6194] = f[303] && f[485] && f[207] && !f[354];
	assign leaf[6195] = f[303] && f[485] && f[207] && f[354];
	
	// Tree 429, Classifier 9, Iteration: 42
	assign leaf[6196] = !f[350] && !f[406] && !f[487] && !f[514];
	assign leaf[6197] = !f[350] && !f[406] && !f[487] && f[514];
	assign leaf[6198] = !f[350] && !f[406] && f[487] && !f[404];
	assign leaf[6199] = !f[350] && !f[406] && f[487] && f[404];
	assign leaf[6200] = !f[350] && f[406] && !f[292] && !f[462];
	assign leaf[6201] = !f[350] && f[406] && !f[292] && f[462];
	assign leaf[6202] = !f[350] && f[406] && f[292] && !f[181];
	assign leaf[6203] = !f[350] && f[406] && f[292] && f[181];
	assign leaf[6204] = f[350] && !f[487] && !f[324] && !f[608];
	assign leaf[6205] = f[350] && !f[487] && !f[324] && f[608];
	assign leaf[6206] = f[350] && !f[487] && f[324] && !f[461];
	assign leaf[6207] = f[350] && !f[487] && f[324] && f[461];
	assign leaf[6208] = f[350] && f[487] && !f[434] && !f[580];
	assign leaf[6209] = f[350] && f[487] && !f[434] && f[580];
	assign leaf[6210] = f[350] && f[487] && f[434] && !f[600];
	assign leaf[6211] = f[350] && f[487] && f[434] && f[600];
	
	// Tree 430, Classifier 0, Iteration: 43
	assign leaf[6212] = !f[408] && !f[491] && !f[209] && !f[150];
	assign leaf[6213] = !f[408] && !f[491] && !f[209] && f[150];
	assign leaf[6214] = !f[408] && !f[491] && f[209] && !f[488];
	assign leaf[6215] = !f[408] && !f[491] && f[209] && f[488];
	assign leaf[6216] = !f[408] && f[491] && !f[210] && !f[576];
	assign leaf[6217] = !f[408] && f[491] && !f[210] && f[576];
	assign leaf[6218] = !f[408] && f[491] && f[210] && !f[410];
	assign leaf[6219] = !f[408] && f[491] && f[210] && f[410];
	assign leaf[6220] = f[408] && !f[268] && !f[427];
	assign leaf[6221] = f[408] && !f[268] && f[427] && !f[595];
	assign leaf[6222] = f[408] && !f[268] && f[427] && f[595];
	assign leaf[6223] = f[408] && f[268] && !f[514] && !f[271];
	assign leaf[6224] = f[408] && f[268] && !f[514] && f[271];
	assign leaf[6225] = f[408] && f[268] && f[514] && !f[656];
	assign leaf[6226] = f[408] && f[268] && f[514] && f[656];
	
	// Tree 431, Classifier 1, Iteration: 43
	assign leaf[6227] = !f[176] && !f[271] && !f[189] && !f[266];
	assign leaf[6228] = !f[176] && !f[271] && !f[189] && f[266];
	assign leaf[6229] = !f[176] && !f[271] && f[189] && !f[491];
	assign leaf[6230] = !f[176] && !f[271] && f[189] && f[491];
	assign leaf[6231] = !f[176] && f[271] && !f[381] && !f[573];
	assign leaf[6232] = !f[176] && f[271] && !f[381] && f[573];
	assign leaf[6233] = !f[176] && f[271] && f[381] && !f[296];
	assign leaf[6234] = !f[176] && f[271] && f[381] && f[296];
	assign leaf[6235] = f[176] && !f[290] && !f[127];
	assign leaf[6236] = f[176] && !f[290] && f[127];
	assign leaf[6237] = f[176] && f[290];
	
	// Tree 432, Classifier 2, Iteration: 43
	assign leaf[6238] = !f[486] && !f[432] && !f[512] && !f[689];
	assign leaf[6239] = !f[486] && !f[432] && !f[512] && f[689];
	assign leaf[6240] = !f[486] && !f[432] && f[512] && !f[404];
	assign leaf[6241] = !f[486] && !f[432] && f[512] && f[404];
	assign leaf[6242] = !f[486] && f[432] && !f[455] && !f[403];
	assign leaf[6243] = !f[486] && f[432] && !f[455] && f[403];
	assign leaf[6244] = !f[486] && f[432] && f[455] && !f[465];
	assign leaf[6245] = !f[486] && f[432] && f[455] && f[465];
	assign leaf[6246] = f[486] && !f[690] && !f[687] && !f[383];
	assign leaf[6247] = f[486] && !f[690] && !f[687] && f[383];
	assign leaf[6248] = f[486] && !f[690] && f[687] && !f[598];
	assign leaf[6249] = f[486] && !f[690] && f[687] && f[598];
	assign leaf[6250] = f[486] && f[690] && !f[657] && !f[573];
	assign leaf[6251] = f[486] && f[690] && !f[657] && f[573];
	assign leaf[6252] = f[486] && f[690] && f[657];
	
	// Tree 433, Classifier 3, Iteration: 43
	assign leaf[6253] = !f[708] && !f[120] && !f[318] && !f[344];
	assign leaf[6254] = !f[708] && !f[120] && !f[318] && f[344];
	assign leaf[6255] = !f[708] && !f[120] && f[318] && !f[293];
	assign leaf[6256] = !f[708] && !f[120] && f[318] && f[293];
	assign leaf[6257] = !f[708] && f[120] && !f[292] && !f[345];
	assign leaf[6258] = !f[708] && f[120] && !f[292] && f[345];
	assign leaf[6259] = !f[708] && f[120] && f[292] && !f[260];
	assign leaf[6260] = !f[708] && f[120] && f[292] && f[260];
	assign leaf[6261] = f[708] && !f[599] && !f[463] && !f[377];
	assign leaf[6262] = f[708] && !f[599] && !f[463] && f[377];
	assign leaf[6263] = f[708] && !f[599] && f[463] && !f[382];
	assign leaf[6264] = f[708] && !f[599] && f[463] && f[382];
	assign leaf[6265] = f[708] && f[599] && !f[602];
	assign leaf[6266] = f[708] && f[599] && f[602];
	
	// Tree 434, Classifier 4, Iteration: 43
	assign leaf[6267] = !f[398] && !f[403] && !f[181] && !f[206];
	assign leaf[6268] = !f[398] && !f[403] && !f[181] && f[206];
	assign leaf[6269] = !f[398] && !f[403] && f[181] && !f[184];
	assign leaf[6270] = !f[398] && !f[403] && f[181] && f[184];
	assign leaf[6271] = !f[398] && f[403] && !f[469] && !f[128];
	assign leaf[6272] = !f[398] && f[403] && !f[469] && f[128];
	assign leaf[6273] = !f[398] && f[403] && f[469] && !f[213];
	assign leaf[6274] = !f[398] && f[403] && f[469] && f[213];
	assign leaf[6275] = f[398] && !f[331] && !f[555] && !f[327];
	assign leaf[6276] = f[398] && !f[331] && !f[555] && f[327];
	assign leaf[6277] = f[398] && !f[331] && f[555] && !f[323];
	assign leaf[6278] = f[398] && !f[331] && f[555] && f[323];
	assign leaf[6279] = f[398] && f[331] && !f[461] && !f[382];
	assign leaf[6280] = f[398] && f[331] && !f[461] && f[382];
	assign leaf[6281] = f[398] && f[331] && f[461] && !f[241];
	assign leaf[6282] = f[398] && f[331] && f[461] && f[241];
	
	// Tree 435, Classifier 5, Iteration: 43
	assign leaf[6283] = !f[488] && !f[485] && !f[133] && !f[380];
	assign leaf[6284] = !f[488] && !f[485] && !f[133] && f[380];
	assign leaf[6285] = !f[488] && !f[485] && f[133] && !f[218];
	assign leaf[6286] = !f[488] && !f[485] && f[133] && f[218];
	assign leaf[6287] = !f[488] && f[485] && !f[430] && !f[372];
	assign leaf[6288] = !f[488] && f[485] && !f[430] && f[372];
	assign leaf[6289] = !f[488] && f[485] && f[430] && !f[541];
	assign leaf[6290] = !f[488] && f[485] && f[430] && f[541];
	assign leaf[6291] = f[488] && !f[717] && !f[430] && !f[183];
	assign leaf[6292] = f[488] && !f[717] && !f[430] && f[183];
	assign leaf[6293] = f[488] && !f[717] && f[430] && !f[322];
	assign leaf[6294] = f[488] && !f[717] && f[430] && f[322];
	assign leaf[6295] = f[488] && f[717] && !f[632];
	assign leaf[6296] = f[488] && f[717] && f[632];
	
	// Tree 436, Classifier 6, Iteration: 43
	assign leaf[6297] = !f[275] && !f[101] && !f[163] && !f[268];
	assign leaf[6298] = !f[275] && !f[101] && !f[163] && f[268];
	assign leaf[6299] = !f[275] && !f[101] && f[163] && !f[355];
	assign leaf[6300] = !f[275] && !f[101] && f[163] && f[355];
	assign leaf[6301] = !f[275] && f[101] && !f[74] && !f[547];
	assign leaf[6302] = !f[275] && f[101] && !f[74] && f[547];
	assign leaf[6303] = !f[275] && f[101] && f[74] && !f[485];
	assign leaf[6304] = !f[275] && f[101] && f[74] && f[485];
	assign leaf[6305] = f[275] && !f[272];
	assign leaf[6306] = f[275] && f[272] && !f[332] && !f[515];
	assign leaf[6307] = f[275] && f[272] && !f[332] && f[515];
	assign leaf[6308] = f[275] && f[272] && f[332];
	
	// Tree 437, Classifier 7, Iteration: 43
	assign leaf[6309] = !f[438] && !f[214] && !f[301] && !f[349];
	assign leaf[6310] = !f[438] && !f[214] && !f[301] && f[349];
	assign leaf[6311] = !f[438] && !f[214] && f[301] && !f[541];
	assign leaf[6312] = !f[438] && !f[214] && f[301] && f[541];
	assign leaf[6313] = !f[438] && f[214] && !f[544] && !f[681];
	assign leaf[6314] = !f[438] && f[214] && !f[544] && f[681];
	assign leaf[6315] = !f[438] && f[214] && f[544] && !f[152];
	assign leaf[6316] = !f[438] && f[214] && f[544] && f[152];
	assign leaf[6317] = f[438] && !f[202] && !f[515] && !f[596];
	assign leaf[6318] = f[438] && !f[202] && !f[515] && f[596];
	assign leaf[6319] = f[438] && !f[202] && f[515] && !f[318];
	assign leaf[6320] = f[438] && !f[202] && f[515] && f[318];
	assign leaf[6321] = f[438] && f[202] && !f[257] && !f[598];
	assign leaf[6322] = f[438] && f[202] && !f[257] && f[598];
	assign leaf[6323] = f[438] && f[202] && f[257] && !f[260];
	assign leaf[6324] = f[438] && f[202] && f[257] && f[260];
	
	// Tree 438, Classifier 8, Iteration: 43
	assign leaf[6325] = !f[542] && !f[512] && !f[544] && !f[510];
	assign leaf[6326] = !f[542] && !f[512] && !f[544] && f[510];
	assign leaf[6327] = !f[542] && !f[512] && f[544] && !f[549];
	assign leaf[6328] = !f[542] && !f[512] && f[544] && f[549];
	assign leaf[6329] = !f[542] && f[512] && !f[322] && !f[403];
	assign leaf[6330] = !f[542] && f[512] && !f[322] && f[403];
	assign leaf[6331] = !f[542] && f[512] && f[322] && !f[540];
	assign leaf[6332] = !f[542] && f[512] && f[322] && f[540];
	assign leaf[6333] = f[542] && !f[511] && !f[544] && !f[518];
	assign leaf[6334] = f[542] && !f[511] && !f[544] && f[518];
	assign leaf[6335] = f[542] && !f[511] && f[544] && !f[296];
	assign leaf[6336] = f[542] && !f[511] && f[544] && f[296];
	assign leaf[6337] = f[542] && f[511] && !f[681] && !f[634];
	assign leaf[6338] = f[542] && f[511] && !f[681] && f[634];
	assign leaf[6339] = f[542] && f[511] && f[681] && !f[491];
	assign leaf[6340] = f[542] && f[511] && f[681] && f[491];
	
	// Tree 439, Classifier 9, Iteration: 43
	assign leaf[6341] = !f[472] && !f[201] && !f[315] && !f[205];
	assign leaf[6342] = !f[472] && !f[201] && !f[315] && f[205];
	assign leaf[6343] = !f[472] && !f[201] && f[315] && !f[317];
	assign leaf[6344] = !f[472] && !f[201] && f[315] && f[317];
	assign leaf[6345] = !f[472] && f[201] && !f[666];
	assign leaf[6346] = !f[472] && f[201] && f[666];
	assign leaf[6347] = f[472];
	
	// Tree 440, Classifier 0, Iteration: 44
	assign leaf[6348] = !f[319] && !f[494] && !f[374] && !f[627];
	assign leaf[6349] = !f[319] && !f[494] && !f[374] && f[627];
	assign leaf[6350] = !f[319] && !f[494] && f[374] && !f[376];
	assign leaf[6351] = !f[319] && !f[494] && f[374] && f[376];
	assign leaf[6352] = !f[319] && f[494] && !f[237] && !f[176];
	assign leaf[6353] = !f[319] && f[494] && !f[237] && f[176];
	assign leaf[6354] = !f[319] && f[494] && f[237] && !f[370];
	assign leaf[6355] = !f[319] && f[494] && f[237] && f[370];
	assign leaf[6356] = f[319] && !f[543] && !f[233] && !f[409];
	assign leaf[6357] = f[319] && !f[543] && !f[233] && f[409];
	assign leaf[6358] = f[319] && !f[543] && f[233] && !f[297];
	assign leaf[6359] = f[319] && !f[543] && f[233] && f[297];
	assign leaf[6360] = f[319] && f[543] && !f[541] && !f[625];
	assign leaf[6361] = f[319] && f[543] && !f[541] && f[625];
	assign leaf[6362] = f[319] && f[543] && f[541] && !f[160];
	assign leaf[6363] = f[319] && f[543] && f[541] && f[160];
	
	// Tree 441, Classifier 1, Iteration: 44
	assign leaf[6364] = !f[608] && !f[260] && !f[661] && !f[292];
	assign leaf[6365] = !f[608] && !f[260] && !f[661] && f[292];
	assign leaf[6366] = !f[608] && !f[260] && f[661] && !f[547];
	assign leaf[6367] = !f[608] && !f[260] && f[661] && f[547];
	assign leaf[6368] = !f[608] && f[260] && !f[154];
	assign leaf[6369] = !f[608] && f[260] && f[154];
	assign leaf[6370] = f[608] && !f[488] && !f[548] && !f[625];
	assign leaf[6371] = f[608] && !f[488] && !f[548] && f[625];
	assign leaf[6372] = f[608] && !f[488] && f[548] && !f[267];
	assign leaf[6373] = f[608] && !f[488] && f[548] && f[267];
	assign leaf[6374] = f[608] && f[488] && !f[318] && !f[379];
	assign leaf[6375] = f[608] && f[488] && !f[318] && f[379];
	assign leaf[6376] = f[608] && f[488] && f[318];
	
	// Tree 442, Classifier 2, Iteration: 44
	assign leaf[6377] = !f[677] && !f[323] && !f[261] && !f[292];
	assign leaf[6378] = !f[677] && !f[323] && !f[261] && f[292];
	assign leaf[6379] = !f[677] && !f[323] && f[261] && !f[652];
	assign leaf[6380] = !f[677] && !f[323] && f[261] && f[652];
	assign leaf[6381] = !f[677] && f[323] && !f[326] && !f[516];
	assign leaf[6382] = !f[677] && f[323] && !f[326] && f[516];
	assign leaf[6383] = !f[677] && f[323] && f[326] && !f[578];
	assign leaf[6384] = !f[677] && f[323] && f[326] && f[578];
	assign leaf[6385] = f[677] && !f[158];
	assign leaf[6386] = f[677] && f[158];
	
	// Tree 443, Classifier 3, Iteration: 44
	assign leaf[6387] = !f[427] && !f[486] && !f[124] && !f[554];
	assign leaf[6388] = !f[427] && !f[486] && !f[124] && f[554];
	assign leaf[6389] = !f[427] && !f[486] && f[124] && !f[207];
	assign leaf[6390] = !f[427] && !f[486] && f[124] && f[207];
	assign leaf[6391] = !f[427] && f[486] && !f[541] && !f[542];
	assign leaf[6392] = !f[427] && f[486] && !f[541] && f[542];
	assign leaf[6393] = !f[427] && f[486] && f[541] && !f[483];
	assign leaf[6394] = !f[427] && f[486] && f[541] && f[483];
	assign leaf[6395] = f[427] && !f[158] && !f[710] && !f[466];
	assign leaf[6396] = f[427] && !f[158] && !f[710] && f[466];
	assign leaf[6397] = f[427] && !f[158] && f[710];
	assign leaf[6398] = f[427] && f[158] && !f[356] && !f[494];
	assign leaf[6399] = f[427] && f[158] && !f[356] && f[494];
	assign leaf[6400] = f[427] && f[158] && f[356] && !f[486];
	assign leaf[6401] = f[427] && f[158] && f[356] && f[486];
	
	// Tree 444, Classifier 4, Iteration: 44
	assign leaf[6402] = !f[102] && !f[97] && !f[714] && !f[381];
	assign leaf[6403] = !f[102] && !f[97] && !f[714] && f[381];
	assign leaf[6404] = !f[102] && !f[97] && f[714] && !f[237];
	assign leaf[6405] = !f[102] && !f[97] && f[714] && f[237];
	assign leaf[6406] = !f[102] && f[97] && !f[573];
	assign leaf[6407] = !f[102] && f[97] && f[573];
	assign leaf[6408] = f[102] && !f[296];
	assign leaf[6409] = f[102] && f[296];
	
	// Tree 445, Classifier 5, Iteration: 44
	assign leaf[6410] = !f[411] && !f[301] && !f[217] && !f[295];
	assign leaf[6411] = !f[411] && !f[301] && !f[217] && f[295];
	assign leaf[6412] = !f[411] && !f[301] && f[217] && !f[298];
	assign leaf[6413] = !f[411] && !f[301] && f[217] && f[298];
	assign leaf[6414] = !f[411] && f[301] && !f[185] && !f[440];
	assign leaf[6415] = !f[411] && f[301] && !f[185] && f[440];
	assign leaf[6416] = !f[411] && f[301] && f[185] && !f[269];
	assign leaf[6417] = !f[411] && f[301] && f[185] && f[269];
	assign leaf[6418] = f[411] && !f[496] && !f[353] && !f[124];
	assign leaf[6419] = f[411] && !f[496] && !f[353] && f[124];
	assign leaf[6420] = f[411] && !f[496] && f[353] && !f[299];
	assign leaf[6421] = f[411] && !f[496] && f[353] && f[299];
	assign leaf[6422] = f[411] && f[496] && !f[185] && !f[127];
	assign leaf[6423] = f[411] && f[496] && !f[185] && f[127];
	assign leaf[6424] = f[411] && f[496] && f[185] && !f[271];
	assign leaf[6425] = f[411] && f[496] && f[185] && f[271];
	
	// Tree 446, Classifier 6, Iteration: 44
	assign leaf[6426] = !f[517] && !f[178] && !f[600] && !f[317];
	assign leaf[6427] = !f[517] && !f[178] && !f[600] && f[317];
	assign leaf[6428] = !f[517] && !f[178] && f[600] && !f[574];
	assign leaf[6429] = !f[517] && !f[178] && f[600] && f[574];
	assign leaf[6430] = !f[517] && f[178] && !f[319] && !f[184];
	assign leaf[6431] = !f[517] && f[178] && !f[319] && f[184];
	assign leaf[6432] = !f[517] && f[178] && f[319] && !f[428];
	assign leaf[6433] = !f[517] && f[178] && f[319] && f[428];
	assign leaf[6434] = f[517] && !f[652] && !f[602] && !f[383];
	assign leaf[6435] = f[517] && !f[652] && !f[602] && f[383];
	assign leaf[6436] = f[517] && !f[652] && f[602] && !f[381];
	assign leaf[6437] = f[517] && !f[652] && f[602] && f[381];
	assign leaf[6438] = f[517] && f[652];
	
	// Tree 447, Classifier 7, Iteration: 44
	assign leaf[6439] = !f[715] && !f[576] && !f[632] && !f[179];
	assign leaf[6440] = !f[715] && !f[576] && !f[632] && f[179];
	assign leaf[6441] = !f[715] && !f[576] && f[632] && !f[716];
	assign leaf[6442] = !f[715] && !f[576] && f[632] && f[716];
	assign leaf[6443] = !f[715] && f[576] && !f[230] && !f[406];
	assign leaf[6444] = !f[715] && f[576] && !f[230] && f[406];
	assign leaf[6445] = !f[715] && f[576] && f[230] && !f[492];
	assign leaf[6446] = !f[715] && f[576] && f[230] && f[492];
	assign leaf[6447] = f[715] && !f[631] && !f[181] && !f[518];
	assign leaf[6448] = f[715] && !f[631] && !f[181] && f[518];
	assign leaf[6449] = f[715] && !f[631] && f[181] && !f[322];
	assign leaf[6450] = f[715] && !f[631] && f[181] && f[322];
	assign leaf[6451] = f[715] && f[631] && !f[518] && !f[436];
	assign leaf[6452] = f[715] && f[631] && !f[518] && f[436];
	assign leaf[6453] = f[715] && f[631] && f[518] && !f[302];
	assign leaf[6454] = f[715] && f[631] && f[518] && f[302];
	
	// Tree 448, Classifier 8, Iteration: 44
	assign leaf[6455] = !f[341] && !f[688] && !f[542] && !f[511];
	assign leaf[6456] = !f[341] && !f[688] && !f[542] && f[511];
	assign leaf[6457] = !f[341] && !f[688] && f[542] && !f[511];
	assign leaf[6458] = !f[341] && !f[688] && f[542] && f[511];
	assign leaf[6459] = !f[341] && f[688] && !f[632] && !f[550];
	assign leaf[6460] = !f[341] && f[688] && !f[632] && f[550];
	assign leaf[6461] = !f[341] && f[688] && f[632] && !f[546];
	assign leaf[6462] = !f[341] && f[688] && f[632] && f[546];
	assign leaf[6463] = f[341] && !f[315] && !f[636];
	assign leaf[6464] = f[341] && !f[315] && f[636];
	assign leaf[6465] = f[341] && f[315] && !f[491] && !f[487];
	assign leaf[6466] = f[341] && f[315] && !f[491] && f[487];
	assign leaf[6467] = f[341] && f[315] && f[491] && !f[350];
	assign leaf[6468] = f[341] && f[315] && f[491] && f[350];
	
	// Tree 449, Classifier 9, Iteration: 44
	assign leaf[6469] = !f[740] && !f[742] && !f[709] && !f[182];
	assign leaf[6470] = !f[740] && !f[742] && !f[709] && f[182];
	assign leaf[6471] = !f[740] && !f[742] && f[709] && !f[236];
	assign leaf[6472] = !f[740] && !f[742] && f[709] && f[236];
	assign leaf[6473] = !f[740] && f[742] && !f[242] && !f[268];
	assign leaf[6474] = !f[740] && f[742] && !f[242] && f[268];
	assign leaf[6475] = !f[740] && f[742] && f[242] && !f[206];
	assign leaf[6476] = !f[740] && f[742] && f[242] && f[206];
	assign leaf[6477] = f[740] && !f[243] && !f[406] && !f[711];
	assign leaf[6478] = f[740] && !f[243] && !f[406] && f[711];
	assign leaf[6479] = f[740] && !f[243] && f[406] && !f[377];
	assign leaf[6480] = f[740] && !f[243] && f[406] && f[377];
	assign leaf[6481] = f[740] && f[243] && !f[235] && !f[404];
	assign leaf[6482] = f[740] && f[243] && !f[235] && f[404];
	assign leaf[6483] = f[740] && f[243] && f[235] && !f[349];
	assign leaf[6484] = f[740] && f[243] && f[235] && f[349];
	
	// Tree 450, Classifier 0, Iteration: 45
	assign leaf[6485] = !f[444] && !f[375] && !f[520] && !f[293];
	assign leaf[6486] = !f[444] && !f[375] && !f[520] && f[293];
	assign leaf[6487] = !f[444] && !f[375] && f[520] && !f[373];
	assign leaf[6488] = !f[444] && !f[375] && f[520] && f[373];
	assign leaf[6489] = !f[444] && f[375] && !f[486] && !f[352];
	assign leaf[6490] = !f[444] && f[375] && !f[486] && f[352];
	assign leaf[6491] = !f[444] && f[375] && f[486] && !f[99];
	assign leaf[6492] = !f[444] && f[375] && f[486] && f[99];
	assign leaf[6493] = f[444] && !f[437] && !f[370];
	assign leaf[6494] = f[444] && !f[437] && f[370] && !f[379];
	assign leaf[6495] = f[444] && !f[437] && f[370] && f[379];
	assign leaf[6496] = f[444] && f[437];
	
	// Tree 451, Classifier 1, Iteration: 45
	assign leaf[6497] = !f[578] && !f[148] && !f[289] && !f[99];
	assign leaf[6498] = !f[578] && !f[148] && !f[289] && f[99];
	assign leaf[6499] = !f[578] && !f[148] && f[289] && !f[627];
	assign leaf[6500] = !f[578] && !f[148] && f[289] && f[627];
	assign leaf[6501] = !f[578] && f[148];
	assign leaf[6502] = f[578] && !f[519] && !f[608] && !f[262];
	assign leaf[6503] = f[578] && !f[519] && !f[608] && f[262];
	assign leaf[6504] = f[578] && !f[519] && f[608] && !f[405];
	assign leaf[6505] = f[578] && !f[519] && f[608] && f[405];
	assign leaf[6506] = f[578] && f[519] && !f[461] && !f[350];
	assign leaf[6507] = f[578] && f[519] && !f[461] && f[350];
	assign leaf[6508] = f[578] && f[519] && f[461] && !f[263];
	assign leaf[6509] = f[578] && f[519] && f[461] && f[263];
	
	// Tree 452, Classifier 2, Iteration: 45
	assign leaf[6510] = !f[681] && !f[461] && !f[573] && !f[430];
	assign leaf[6511] = !f[681] && !f[461] && !f[573] && f[430];
	assign leaf[6512] = !f[681] && !f[461] && f[573] && !f[204];
	assign leaf[6513] = !f[681] && !f[461] && f[573] && f[204];
	assign leaf[6514] = !f[681] && f[461] && !f[525] && !f[388];
	assign leaf[6515] = !f[681] && f[461] && !f[525] && f[388];
	assign leaf[6516] = !f[681] && f[461] && f[525] && !f[607];
	assign leaf[6517] = !f[681] && f[461] && f[525] && f[607];
	assign leaf[6518] = f[681] && !f[603] && !f[686] && !f[462];
	assign leaf[6519] = f[681] && !f[603] && !f[686] && f[462];
	assign leaf[6520] = f[681] && !f[603] && f[686] && !f[631];
	assign leaf[6521] = f[681] && !f[603] && f[686] && f[631];
	assign leaf[6522] = f[681] && f[603] && !f[432] && !f[685];
	assign leaf[6523] = f[681] && f[603] && !f[432] && f[685];
	assign leaf[6524] = f[681] && f[603] && f[432] && !f[594];
	assign leaf[6525] = f[681] && f[603] && f[432] && f[594];
	
	// Tree 453, Classifier 3, Iteration: 45
	assign leaf[6526] = !f[451] && !f[133] && !f[591] && !f[210];
	assign leaf[6527] = !f[451] && !f[133] && !f[591] && f[210];
	assign leaf[6528] = !f[451] && !f[133] && f[591] && !f[404];
	assign leaf[6529] = !f[451] && !f[133] && f[591] && f[404];
	assign leaf[6530] = !f[451] && f[133] && !f[272] && !f[179];
	assign leaf[6531] = !f[451] && f[133] && !f[272] && f[179];
	assign leaf[6532] = !f[451] && f[133] && f[272] && !f[462];
	assign leaf[6533] = !f[451] && f[133] && f[272] && f[462];
	assign leaf[6534] = f[451] && !f[352];
	assign leaf[6535] = f[451] && f[352] && !f[159];
	assign leaf[6536] = f[451] && f[352] && f[159];
	
	// Tree 454, Classifier 4, Iteration: 45
	assign leaf[6537] = !f[179] && !f[635] && !f[241] && !f[158];
	assign leaf[6538] = !f[179] && !f[635] && !f[241] && f[158];
	assign leaf[6539] = !f[179] && !f[635] && f[241] && !f[244];
	assign leaf[6540] = !f[179] && !f[635] && f[241] && f[244];
	assign leaf[6541] = !f[179] && f[635] && !f[747] && !f[660];
	assign leaf[6542] = !f[179] && f[635] && !f[747] && f[660];
	assign leaf[6543] = !f[179] && f[635] && f[747];
	assign leaf[6544] = f[179] && !f[181] && !f[204] && !f[153];
	assign leaf[6545] = f[179] && !f[181] && !f[204] && f[153];
	assign leaf[6546] = f[179] && !f[181] && f[204] && !f[300];
	assign leaf[6547] = f[179] && !f[181] && f[204] && f[300];
	assign leaf[6548] = f[179] && f[181] && !f[263] && !f[273];
	assign leaf[6549] = f[179] && f[181] && !f[263] && f[273];
	assign leaf[6550] = f[179] && f[181] && f[263] && !f[183];
	assign leaf[6551] = f[179] && f[181] && f[263] && f[183];
	
	// Tree 455, Classifier 5, Iteration: 45
	assign leaf[6552] = !f[556] && !f[654] && !f[459] && !f[543];
	assign leaf[6553] = !f[556] && !f[654] && !f[459] && f[543];
	assign leaf[6554] = !f[556] && !f[654] && f[459] && !f[401];
	assign leaf[6555] = !f[556] && !f[654] && f[459] && f[401];
	assign leaf[6556] = !f[556] && f[654] && !f[264] && !f[153];
	assign leaf[6557] = !f[556] && f[654] && !f[264] && f[153];
	assign leaf[6558] = !f[556] && f[654] && f[264] && !f[320];
	assign leaf[6559] = !f[556] && f[654] && f[264] && f[320];
	assign leaf[6560] = f[556] && !f[372];
	assign leaf[6561] = f[556] && f[372] && !f[526];
	assign leaf[6562] = f[556] && f[372] && f[526] && !f[636];
	assign leaf[6563] = f[556] && f[372] && f[526] && f[636];
	
	// Tree 456, Classifier 6, Iteration: 45
	assign leaf[6564] = !f[682] && !f[459] && !f[387] && !f[429];
	assign leaf[6565] = !f[682] && !f[459] && !f[387] && f[429];
	assign leaf[6566] = !f[682] && !f[459] && f[387] && !f[409];
	assign leaf[6567] = !f[682] && !f[459] && f[387] && f[409];
	assign leaf[6568] = !f[682] && f[459] && !f[544] && !f[159];
	assign leaf[6569] = !f[682] && f[459] && !f[544] && f[159];
	assign leaf[6570] = !f[682] && f[459] && f[544] && !f[487];
	assign leaf[6571] = !f[682] && f[459] && f[544] && f[487];
	assign leaf[6572] = f[682];
	
	// Tree 457, Classifier 7, Iteration: 45
	assign leaf[6573] = !f[128] && !f[241] && !f[322] && !f[434];
	assign leaf[6574] = !f[128] && !f[241] && !f[322] && f[434];
	assign leaf[6575] = !f[128] && !f[241] && f[322] && !f[412];
	assign leaf[6576] = !f[128] && !f[241] && f[322] && f[412];
	assign leaf[6577] = !f[128] && f[241] && !f[239] && !f[154];
	assign leaf[6578] = !f[128] && f[241] && !f[239] && f[154];
	assign leaf[6579] = !f[128] && f[241] && f[239] && !f[207];
	assign leaf[6580] = !f[128] && f[241] && f[239] && f[207];
	assign leaf[6581] = f[128];
	
	// Tree 458, Classifier 8, Iteration: 45
	assign leaf[6582] = !f[325] && !f[354] && !f[268] && !f[356];
	assign leaf[6583] = !f[325] && !f[354] && !f[268] && f[356];
	assign leaf[6584] = !f[325] && !f[354] && f[268] && !f[632];
	assign leaf[6585] = !f[325] && !f[354] && f[268] && f[632];
	assign leaf[6586] = !f[325] && f[354] && !f[411] && !f[593];
	assign leaf[6587] = !f[325] && f[354] && !f[411] && f[593];
	assign leaf[6588] = !f[325] && f[354] && f[411] && !f[554];
	assign leaf[6589] = !f[325] && f[354] && f[411] && f[554];
	assign leaf[6590] = f[325] && !f[409] && !f[492] && !f[518];
	assign leaf[6591] = f[325] && !f[409] && !f[492] && f[518];
	assign leaf[6592] = f[325] && !f[409] && f[492] && !f[403];
	assign leaf[6593] = f[325] && !f[409] && f[492] && f[403];
	assign leaf[6594] = f[325] && f[409] && !f[495] && !f[351];
	assign leaf[6595] = f[325] && f[409] && !f[495] && f[351];
	assign leaf[6596] = f[325] && f[409] && f[495] && !f[426];
	assign leaf[6597] = f[325] && f[409] && f[495] && f[426];
	
	// Tree 459, Classifier 9, Iteration: 45
	assign leaf[6598] = !f[746] && !f[734] && !f[275] && !f[606];
	assign leaf[6599] = !f[746] && !f[734] && !f[275] && f[606];
	assign leaf[6600] = !f[746] && !f[734] && f[275] && !f[215];
	assign leaf[6601] = !f[746] && !f[734] && f[275] && f[215];
	assign leaf[6602] = !f[746] && f[734] && !f[431];
	assign leaf[6603] = !f[746] && f[734] && f[431];
	assign leaf[6604] = f[746] && !f[431] && !f[291] && !f[243];
	assign leaf[6605] = f[746] && !f[431] && !f[291] && f[243];
	assign leaf[6606] = f[746] && !f[431] && f[291] && !f[401];
	assign leaf[6607] = f[746] && !f[431] && f[291] && f[401];
	assign leaf[6608] = f[746] && f[431] && !f[661];
	assign leaf[6609] = f[746] && f[431] && f[661];
	
	// Tree 460, Classifier 0, Iteration: 46
	assign leaf[6610] = !f[434] && !f[664] && !f[379] && !f[332];
	assign leaf[6611] = !f[434] && !f[664] && !f[379] && f[332];
	assign leaf[6612] = !f[434] && !f[664] && f[379] && !f[488];
	assign leaf[6613] = !f[434] && !f[664] && f[379] && f[488];
	assign leaf[6614] = !f[434] && f[664] && !f[178];
	assign leaf[6615] = !f[434] && f[664] && f[178] && !f[498];
	assign leaf[6616] = !f[434] && f[664] && f[178] && f[498];
	assign leaf[6617] = f[434] && !f[436] && !f[185];
	assign leaf[6618] = f[434] && !f[436] && f[185] && !f[457];
	assign leaf[6619] = f[434] && !f[436] && f[185] && f[457];
	assign leaf[6620] = f[434] && f[436] && !f[433] && !f[595];
	assign leaf[6621] = f[434] && f[436] && !f[433] && f[595];
	assign leaf[6622] = f[434] && f[436] && f[433] && !f[414];
	assign leaf[6623] = f[434] && f[436] && f[433] && f[414];
	
	// Tree 461, Classifier 1, Iteration: 46
	assign leaf[6624] = !f[578] && !f[148] && !f[493] && !f[320];
	assign leaf[6625] = !f[578] && !f[148] && !f[493] && f[320];
	assign leaf[6626] = !f[578] && !f[148] && f[493] && !f[237];
	assign leaf[6627] = !f[578] && !f[148] && f[493] && f[237];
	assign leaf[6628] = !f[578] && f[148];
	assign leaf[6629] = f[578] && !f[460] && !f[491] && !f[570];
	assign leaf[6630] = f[578] && !f[460] && !f[491] && f[570];
	assign leaf[6631] = f[578] && !f[460] && f[491] && !f[595];
	assign leaf[6632] = f[578] && !f[460] && f[491] && f[595];
	assign leaf[6633] = f[578] && f[460] && !f[319] && !f[487];
	assign leaf[6634] = f[578] && f[460] && !f[319] && f[487];
	assign leaf[6635] = f[578] && f[460] && f[319] && !f[213];
	assign leaf[6636] = f[578] && f[460] && f[319] && f[213];
	
	// Tree 462, Classifier 2, Iteration: 46
	assign leaf[6637] = !f[324] && !f[509] && !f[571] && !f[267];
	assign leaf[6638] = !f[324] && !f[509] && !f[571] && f[267];
	assign leaf[6639] = !f[324] && !f[509] && f[571] && !f[297];
	assign leaf[6640] = !f[324] && !f[509] && f[571] && f[297];
	assign leaf[6641] = !f[324] && f[509] && !f[457] && !f[403];
	assign leaf[6642] = !f[324] && f[509] && !f[457] && f[403];
	assign leaf[6643] = !f[324] && f[509] && f[457] && !f[376];
	assign leaf[6644] = !f[324] && f[509] && f[457] && f[376];
	assign leaf[6645] = f[324] && !f[347] && !f[356] && !f[215];
	assign leaf[6646] = f[324] && !f[347] && !f[356] && f[215];
	assign leaf[6647] = f[324] && !f[347] && f[356] && !f[204];
	assign leaf[6648] = f[324] && !f[347] && f[356] && f[204];
	assign leaf[6649] = f[324] && f[347] && !f[96] && !f[453];
	assign leaf[6650] = f[324] && f[347] && !f[96] && f[453];
	assign leaf[6651] = f[324] && f[347] && f[96];
	
	// Tree 463, Classifier 3, Iteration: 46
	assign leaf[6652] = !f[458] && !f[566] && !f[266] && !f[355];
	assign leaf[6653] = !f[458] && !f[566] && !f[266] && f[355];
	assign leaf[6654] = !f[458] && !f[566] && f[266] && !f[468];
	assign leaf[6655] = !f[458] && !f[566] && f[266] && f[468];
	assign leaf[6656] = !f[458] && f[566] && !f[517] && !f[455];
	assign leaf[6657] = !f[458] && f[566] && !f[517] && f[455];
	assign leaf[6658] = !f[458] && f[566] && f[517] && !f[621];
	assign leaf[6659] = !f[458] && f[566] && f[517] && f[621];
	assign leaf[6660] = f[458] && !f[489] && !f[540] && !f[653];
	assign leaf[6661] = f[458] && !f[489] && !f[540] && f[653];
	assign leaf[6662] = f[458] && !f[489] && f[540] && !f[372];
	assign leaf[6663] = f[458] && !f[489] && f[540] && f[372];
	assign leaf[6664] = f[458] && f[489] && !f[605] && !f[436];
	assign leaf[6665] = f[458] && f[489] && !f[605] && f[436];
	assign leaf[6666] = f[458] && f[489] && f[605] && !f[346];
	assign leaf[6667] = f[458] && f[489] && f[605] && f[346];
	
	// Tree 464, Classifier 4, Iteration: 46
	assign leaf[6668] = !f[220] && !f[163] && !f[301] && !f[490];
	assign leaf[6669] = !f[220] && !f[163] && !f[301] && f[490];
	assign leaf[6670] = !f[220] && !f[163] && f[301] && !f[384];
	assign leaf[6671] = !f[220] && !f[163] && f[301] && f[384];
	assign leaf[6672] = !f[220] && f[163] && !f[187] && !f[596];
	assign leaf[6673] = !f[220] && f[163] && !f[187] && f[596];
	assign leaf[6674] = !f[220] && f[163] && f[187];
	assign leaf[6675] = f[220] && !f[214] && !f[210] && !f[464];
	assign leaf[6676] = f[220] && !f[214] && !f[210] && f[464];
	assign leaf[6677] = f[220] && !f[214] && f[210] && !f[191];
	assign leaf[6678] = f[220] && !f[214] && f[210] && f[191];
	assign leaf[6679] = f[220] && f[214];
	
	// Tree 465, Classifier 5, Iteration: 46
	assign leaf[6680] = !f[433] && !f[347] && !f[293] && !f[547];
	assign leaf[6681] = !f[433] && !f[347] && !f[293] && f[547];
	assign leaf[6682] = !f[433] && !f[347] && f[293] && !f[258];
	assign leaf[6683] = !f[433] && !f[347] && f[293] && f[258];
	assign leaf[6684] = !f[433] && f[347] && !f[315] && !f[175];
	assign leaf[6685] = !f[433] && f[347] && !f[315] && f[175];
	assign leaf[6686] = !f[433] && f[347] && f[315] && !f[483];
	assign leaf[6687] = !f[433] && f[347] && f[315] && f[483];
	assign leaf[6688] = f[433] && !f[352] && !f[382] && !f[385];
	assign leaf[6689] = f[433] && !f[352] && !f[382] && f[385];
	assign leaf[6690] = f[433] && !f[352] && f[382] && !f[606];
	assign leaf[6691] = f[433] && !f[352] && f[382] && f[606];
	assign leaf[6692] = f[433] && f[352] && !f[331] && !f[468];
	assign leaf[6693] = f[433] && f[352] && !f[331] && f[468];
	assign leaf[6694] = f[433] && f[352] && f[331] && !f[275];
	assign leaf[6695] = f[433] && f[352] && f[331] && f[275];
	
	// Tree 466, Classifier 6, Iteration: 46
	assign leaf[6696] = !f[622] && !f[132] && !f[267] && !f[213];
	assign leaf[6697] = !f[622] && !f[132] && !f[267] && f[213];
	assign leaf[6698] = !f[622] && !f[132] && f[267] && !f[263];
	assign leaf[6699] = !f[622] && !f[132] && f[267] && f[263];
	assign leaf[6700] = !f[622] && f[132] && !f[326] && !f[233];
	assign leaf[6701] = !f[622] && f[132] && !f[326] && f[233];
	assign leaf[6702] = !f[622] && f[132] && f[326] && !f[496];
	assign leaf[6703] = !f[622] && f[132] && f[326] && f[496];
	assign leaf[6704] = f[622];
	
	// Tree 467, Classifier 7, Iteration: 46
	assign leaf[6705] = !f[256] && !f[663] && !f[177] && !f[232];
	assign leaf[6706] = !f[256] && !f[663] && !f[177] && f[232];
	assign leaf[6707] = !f[256] && !f[663] && f[177] && !f[183];
	assign leaf[6708] = !f[256] && !f[663] && f[177] && f[183];
	assign leaf[6709] = !f[256] && f[663] && !f[263] && !f[550];
	assign leaf[6710] = !f[256] && f[663] && !f[263] && f[550];
	assign leaf[6711] = !f[256] && f[663] && f[263] && !f[459];
	assign leaf[6712] = !f[256] && f[663] && f[263] && f[459];
	assign leaf[6713] = f[256] && !f[493] && !f[436];
	assign leaf[6714] = f[256] && !f[493] && f[436] && !f[239];
	assign leaf[6715] = f[256] && !f[493] && f[436] && f[239];
	assign leaf[6716] = f[256] && f[493] && !f[581] && !f[552];
	assign leaf[6717] = f[256] && f[493] && !f[581] && f[552];
	assign leaf[6718] = f[256] && f[493] && f[581];
	
	// Tree 468, Classifier 8, Iteration: 46
	assign leaf[6719] = !f[649] && !f[201] && !f[663] && !f[494];
	assign leaf[6720] = !f[649] && !f[201] && !f[663] && f[494];
	assign leaf[6721] = !f[649] && !f[201] && f[663] && !f[574];
	assign leaf[6722] = !f[649] && !f[201] && f[663] && f[574];
	assign leaf[6723] = !f[649] && f[201] && !f[318] && !f[342];
	assign leaf[6724] = !f[649] && f[201] && !f[318] && f[342];
	assign leaf[6725] = !f[649] && f[201] && f[318] && !f[296];
	assign leaf[6726] = !f[649] && f[201] && f[318] && f[296];
	assign leaf[6727] = f[649] && !f[624] && !f[568];
	assign leaf[6728] = f[649] && !f[624] && f[568];
	assign leaf[6729] = f[649] && f[624] && !f[456] && !f[348];
	assign leaf[6730] = f[649] && f[624] && !f[456] && f[348];
	assign leaf[6731] = f[649] && f[624] && f[456] && !f[437];
	assign leaf[6732] = f[649] && f[624] && f[456] && f[437];
	
	// Tree 469, Classifier 9, Iteration: 46
	assign leaf[6733] = !f[368] && !f[415] && !f[353] && !f[405];
	assign leaf[6734] = !f[368] && !f[415] && !f[353] && f[405];
	assign leaf[6735] = !f[368] && !f[415] && f[353] && !f[378];
	assign leaf[6736] = !f[368] && !f[415] && f[353] && f[378];
	assign leaf[6737] = !f[368] && f[415] && !f[313] && !f[682];
	assign leaf[6738] = !f[368] && f[415] && !f[313] && f[682];
	assign leaf[6739] = !f[368] && f[415] && f[313];
	assign leaf[6740] = f[368] && !f[373] && !f[660] && !f[326];
	assign leaf[6741] = f[368] && !f[373] && !f[660] && f[326];
	assign leaf[6742] = f[368] && !f[373] && f[660] && !f[434];
	assign leaf[6743] = f[368] && !f[373] && f[660] && f[434];
	assign leaf[6744] = f[368] && f[373] && !f[286];
	assign leaf[6745] = f[368] && f[373] && f[286] && !f[238];
	assign leaf[6746] = f[368] && f[373] && f[286] && f[238];
	
	// Tree 470, Classifier 0, Iteration: 47
	assign leaf[6747] = !f[714] && !f[710] && !f[427] && !f[431];
	assign leaf[6748] = !f[714] && !f[710] && !f[427] && f[431];
	assign leaf[6749] = !f[714] && !f[710] && f[427] && !f[377];
	assign leaf[6750] = !f[714] && !f[710] && f[427] && f[377];
	assign leaf[6751] = !f[714] && f[710];
	assign leaf[6752] = f[714] && !f[576];
	assign leaf[6753] = f[714] && f[576];
	
	// Tree 471, Classifier 1, Iteration: 47
	assign leaf[6754] = !f[606] && !f[204] && !f[555] && !f[544];
	assign leaf[6755] = !f[606] && !f[204] && !f[555] && f[544];
	assign leaf[6756] = !f[606] && !f[204] && f[555];
	assign leaf[6757] = !f[606] && f[204] && !f[570];
	assign leaf[6758] = !f[606] && f[204] && f[570];
	assign leaf[6759] = f[606] && !f[515] && !f[547] && !f[153];
	assign leaf[6760] = f[606] && !f[515] && !f[547] && f[153];
	assign leaf[6761] = f[606] && !f[515] && f[547] && !f[688];
	assign leaf[6762] = f[606] && !f[515] && f[547] && f[688];
	assign leaf[6763] = f[606] && f[515] && !f[494] && !f[431];
	assign leaf[6764] = f[606] && f[515] && !f[494] && f[431];
	assign leaf[6765] = f[606] && f[515] && f[494] && !f[241];
	assign leaf[6766] = f[606] && f[515] && f[494] && f[241];
	
	// Tree 472, Classifier 2, Iteration: 47
	assign leaf[6767] = !f[367] && !f[665] && !f[219] && !f[104];
	assign leaf[6768] = !f[367] && !f[665] && !f[219] && f[104];
	assign leaf[6769] = !f[367] && !f[665] && f[219] && !f[159];
	assign leaf[6770] = !f[367] && !f[665] && f[219] && f[159];
	assign leaf[6771] = !f[367] && f[665] && !f[553] && !f[551];
	assign leaf[6772] = !f[367] && f[665] && !f[553] && f[551];
	assign leaf[6773] = !f[367] && f[665] && f[553] && !f[546];
	assign leaf[6774] = !f[367] && f[665] && f[553] && f[546];
	assign leaf[6775] = f[367];
	
	// Tree 473, Classifier 3, Iteration: 47
	assign leaf[6776] = !f[712] && !f[377] && !f[537] && !f[571];
	assign leaf[6777] = !f[712] && !f[377] && !f[537] && f[571];
	assign leaf[6778] = !f[712] && !f[377] && f[537] && !f[209];
	assign leaf[6779] = !f[712] && !f[377] && f[537] && f[209];
	assign leaf[6780] = !f[712] && f[377] && !f[484] && !f[318];
	assign leaf[6781] = !f[712] && f[377] && !f[484] && f[318];
	assign leaf[6782] = !f[712] && f[377] && f[484] && !f[515];
	assign leaf[6783] = !f[712] && f[377] && f[484] && f[515];
	assign leaf[6784] = f[712] && !f[600] && !f[319] && !f[345];
	assign leaf[6785] = f[712] && !f[600] && !f[319] && f[345];
	assign leaf[6786] = f[712] && !f[600] && f[319] && !f[348];
	assign leaf[6787] = f[712] && !f[600] && f[319] && f[348];
	assign leaf[6788] = f[712] && f[600] && !f[317];
	assign leaf[6789] = f[712] && f[600] && f[317];
	
	// Tree 474, Classifier 4, Iteration: 47
	assign leaf[6790] = !f[744] && !f[128] && !f[404] && !f[483];
	assign leaf[6791] = !f[744] && !f[128] && !f[404] && f[483];
	assign leaf[6792] = !f[744] && !f[128] && f[404] && !f[496];
	assign leaf[6793] = !f[744] && !f[128] && f[404] && f[496];
	assign leaf[6794] = !f[744] && f[128] && !f[497] && !f[239];
	assign leaf[6795] = !f[744] && f[128] && !f[497] && f[239];
	assign leaf[6796] = !f[744] && f[128] && f[497] && !f[520];
	assign leaf[6797] = !f[744] && f[128] && f[497] && f[520];
	assign leaf[6798] = f[744] && !f[605];
	assign leaf[6799] = f[744] && f[605];
	
	// Tree 475, Classifier 5, Iteration: 47
	assign leaf[6800] = !f[517] && !f[262] && !f[551] && !f[571];
	assign leaf[6801] = !f[517] && !f[262] && !f[551] && f[571];
	assign leaf[6802] = !f[517] && !f[262] && f[551] && !f[236];
	assign leaf[6803] = !f[517] && !f[262] && f[551] && f[236];
	assign leaf[6804] = !f[517] && f[262] && !f[178] && !f[351];
	assign leaf[6805] = !f[517] && f[262] && !f[178] && f[351];
	assign leaf[6806] = !f[517] && f[262] && f[178] && !f[547];
	assign leaf[6807] = !f[517] && f[262] && f[178] && f[547];
	assign leaf[6808] = f[517] && !f[467] && !f[381] && !f[184];
	assign leaf[6809] = f[517] && !f[467] && !f[381] && f[184];
	assign leaf[6810] = f[517] && !f[467] && f[381] && !f[513];
	assign leaf[6811] = f[517] && !f[467] && f[381] && f[513];
	assign leaf[6812] = f[517] && f[467] && !f[540] && !f[663];
	assign leaf[6813] = f[517] && f[467] && !f[540] && f[663];
	assign leaf[6814] = f[517] && f[467] && f[540] && !f[381];
	assign leaf[6815] = f[517] && f[467] && f[540] && f[381];
	
	// Tree 476, Classifier 6, Iteration: 47
	assign leaf[6816] = !f[455] && !f[596] && !f[607] && !f[661];
	assign leaf[6817] = !f[455] && !f[596] && !f[607] && f[661];
	assign leaf[6818] = !f[455] && !f[596] && f[607] && !f[457];
	assign leaf[6819] = !f[455] && !f[596] && f[607] && f[457];
	assign leaf[6820] = !f[455] && f[596] && !f[370] && !f[457];
	assign leaf[6821] = !f[455] && f[596] && !f[370] && f[457];
	assign leaf[6822] = !f[455] && f[596] && f[370];
	assign leaf[6823] = f[455] && !f[601] && !f[275] && !f[546];
	assign leaf[6824] = f[455] && !f[601] && !f[275] && f[546];
	assign leaf[6825] = f[455] && !f[601] && f[275];
	assign leaf[6826] = f[455] && f[601] && !f[186] && !f[238];
	assign leaf[6827] = f[455] && f[601] && !f[186] && f[238];
	assign leaf[6828] = f[455] && f[601] && f[186] && !f[346];
	assign leaf[6829] = f[455] && f[601] && f[186] && f[346];
	
	// Tree 477, Classifier 7, Iteration: 47
	assign leaf[6830] = !f[295] && !f[350] && !f[213] && !f[435];
	assign leaf[6831] = !f[295] && !f[350] && !f[213] && f[435];
	assign leaf[6832] = !f[295] && !f[350] && f[213] && !f[461];
	assign leaf[6833] = !f[295] && !f[350] && f[213] && f[461];
	assign leaf[6834] = !f[295] && f[350] && !f[210] && !f[266];
	assign leaf[6835] = !f[295] && f[350] && !f[210] && f[266];
	assign leaf[6836] = !f[295] && f[350] && f[210] && !f[460];
	assign leaf[6837] = !f[295] && f[350] && f[210] && f[460];
	assign leaf[6838] = f[295] && !f[404] && !f[491] && !f[212];
	assign leaf[6839] = f[295] && !f[404] && !f[491] && f[212];
	assign leaf[6840] = f[295] && !f[404] && f[491] && !f[658];
	assign leaf[6841] = f[295] && !f[404] && f[491] && f[658];
	assign leaf[6842] = f[295] && f[404] && !f[345] && !f[569];
	assign leaf[6843] = f[295] && f[404] && !f[345] && f[569];
	assign leaf[6844] = f[295] && f[404] && f[345] && !f[406];
	assign leaf[6845] = f[295] && f[404] && f[345] && f[406];
	
	// Tree 478, Classifier 8, Iteration: 47
	assign leaf[6846] = !f[238] && !f[321] && !f[347] && !f[374];
	assign leaf[6847] = !f[238] && !f[321] && !f[347] && f[374];
	assign leaf[6848] = !f[238] && !f[321] && f[347] && !f[402];
	assign leaf[6849] = !f[238] && !f[321] && f[347] && f[402];
	assign leaf[6850] = !f[238] && f[321] && !f[346] && !f[154];
	assign leaf[6851] = !f[238] && f[321] && !f[346] && f[154];
	assign leaf[6852] = !f[238] && f[321] && f[346] && !f[456];
	assign leaf[6853] = !f[238] && f[321] && f[346] && f[456];
	assign leaf[6854] = f[238] && !f[304] && !f[188] && !f[663];
	assign leaf[6855] = f[238] && !f[304] && !f[188] && f[663];
	assign leaf[6856] = f[238] && !f[304] && f[188] && !f[633];
	assign leaf[6857] = f[238] && !f[304] && f[188] && f[633];
	assign leaf[6858] = f[238] && f[304] && !f[400] && !f[520];
	assign leaf[6859] = f[238] && f[304] && !f[400] && f[520];
	assign leaf[6860] = f[238] && f[304] && f[400] && !f[348];
	assign leaf[6861] = f[238] && f[304] && f[400] && f[348];
	
	// Tree 479, Classifier 9, Iteration: 47
	assign leaf[6862] = !f[274] && !f[356] && !f[323] && !f[523];
	assign leaf[6863] = !f[274] && !f[356] && !f[323] && f[523];
	assign leaf[6864] = !f[274] && !f[356] && f[323] && !f[434];
	assign leaf[6865] = !f[274] && !f[356] && f[323] && f[434];
	assign leaf[6866] = !f[274] && f[356] && !f[466] && !f[328];
	assign leaf[6867] = !f[274] && f[356] && !f[466] && f[328];
	assign leaf[6868] = !f[274] && f[356] && f[466] && !f[128];
	assign leaf[6869] = !f[274] && f[356] && f[466] && f[128];
	assign leaf[6870] = f[274] && !f[215] && !f[242] && !f[158];
	assign leaf[6871] = f[274] && !f[215] && !f[242] && f[158];
	assign leaf[6872] = f[274] && !f[215] && f[242] && !f[375];
	assign leaf[6873] = f[274] && !f[215] && f[242] && f[375];
	assign leaf[6874] = f[274] && f[215] && !f[211] && !f[408];
	assign leaf[6875] = f[274] && f[215] && !f[211] && f[408];
	assign leaf[6876] = f[274] && f[215] && f[211] && !f[412];
	assign leaf[6877] = f[274] && f[215] && f[211] && f[412];
	
	// Tree 480, Classifier 0, Iteration: 48
	assign leaf[6878] = !f[238] && !f[219] && !f[266] && !f[464];
	assign leaf[6879] = !f[238] && !f[219] && !f[266] && f[464];
	assign leaf[6880] = !f[238] && !f[219] && f[266] && !f[602];
	assign leaf[6881] = !f[238] && !f[219] && f[266] && f[602];
	assign leaf[6882] = !f[238] && f[219] && !f[510] && !f[189];
	assign leaf[6883] = !f[238] && f[219] && !f[510] && f[189];
	assign leaf[6884] = !f[238] && f[219] && f[510] && !f[241];
	assign leaf[6885] = !f[238] && f[219] && f[510] && f[241];
	assign leaf[6886] = f[238] && !f[269] && !f[625] && !f[386];
	assign leaf[6887] = f[238] && !f[269] && !f[625] && f[386];
	assign leaf[6888] = f[238] && !f[269] && f[625] && !f[325];
	assign leaf[6889] = f[238] && !f[269] && f[625] && f[325];
	assign leaf[6890] = f[238] && f[269] && !f[244] && !f[515];
	assign leaf[6891] = f[238] && f[269] && !f[244] && f[515];
	assign leaf[6892] = f[238] && f[269] && f[244] && !f[295];
	assign leaf[6893] = f[238] && f[269] && f[244] && f[295];
	
	// Tree 481, Classifier 1, Iteration: 48
	assign leaf[6894] = !f[271] && !f[382] && !f[459] && !f[577];
	assign leaf[6895] = !f[271] && !f[382] && !f[459] && f[577];
	assign leaf[6896] = !f[271] && !f[382] && f[459] && !f[377];
	assign leaf[6897] = !f[271] && !f[382] && f[459] && f[377];
	assign leaf[6898] = !f[271] && f[382] && !f[606] && !f[323];
	assign leaf[6899] = !f[271] && f[382] && !f[606] && f[323];
	assign leaf[6900] = !f[271] && f[382] && f[606];
	assign leaf[6901] = f[271] && !f[408] && !f[518] && !f[157];
	assign leaf[6902] = f[271] && !f[408] && !f[518] && f[157];
	assign leaf[6903] = f[271] && !f[408] && f[518];
	assign leaf[6904] = f[271] && f[408] && !f[132] && !f[487];
	assign leaf[6905] = f[271] && f[408] && !f[132] && f[487];
	assign leaf[6906] = f[271] && f[408] && f[132] && !f[156];
	assign leaf[6907] = f[271] && f[408] && f[132] && f[156];
	
	// Tree 482, Classifier 2, Iteration: 48
	assign leaf[6908] = !f[418] && !f[473] && !f[571] && !f[510];
	assign leaf[6909] = !f[418] && !f[473] && !f[571] && f[510];
	assign leaf[6910] = !f[418] && !f[473] && f[571] && !f[715];
	assign leaf[6911] = !f[418] && !f[473] && f[571] && f[715];
	assign leaf[6912] = !f[418] && f[473] && !f[416] && !f[519];
	assign leaf[6913] = !f[418] && f[473] && !f[416] && f[519];
	assign leaf[6914] = !f[418] && f[473] && f[416];
	assign leaf[6915] = f[418];
	
	// Tree 483, Classifier 3, Iteration: 48
	assign leaf[6916] = !f[161] && !f[655] && !f[464] && !f[548];
	assign leaf[6917] = !f[161] && !f[655] && !f[464] && f[548];
	assign leaf[6918] = !f[161] && !f[655] && f[464] && !f[547];
	assign leaf[6919] = !f[161] && !f[655] && f[464] && f[547];
	assign leaf[6920] = !f[161] && f[655] && !f[630] && !f[544];
	assign leaf[6921] = !f[161] && f[655] && !f[630] && f[544];
	assign leaf[6922] = !f[161] && f[655] && f[630] && !f[710];
	assign leaf[6923] = !f[161] && f[655] && f[630] && f[710];
	assign leaf[6924] = f[161] && !f[272] && !f[301] && !f[243];
	assign leaf[6925] = f[161] && !f[272] && !f[301] && f[243];
	assign leaf[6926] = f[161] && !f[272] && f[301];
	assign leaf[6927] = f[161] && f[272] && !f[326] && !f[267];
	assign leaf[6928] = f[161] && f[272] && !f[326] && f[267];
	assign leaf[6929] = f[161] && f[272] && f[326] && !f[460];
	assign leaf[6930] = f[161] && f[272] && f[326] && f[460];
	
	// Tree 484, Classifier 4, Iteration: 48
	assign leaf[6931] = !f[96] && !f[740] && !f[408] && !f[485];
	assign leaf[6932] = !f[96] && !f[740] && !f[408] && f[485];
	assign leaf[6933] = !f[96] && !f[740] && f[408] && !f[348];
	assign leaf[6934] = !f[96] && !f[740] && f[408] && f[348];
	assign leaf[6935] = !f[96] && f[740] && !f[234];
	assign leaf[6936] = !f[96] && f[740] && f[234];
	assign leaf[6937] = f[96] && !f[545];
	assign leaf[6938] = f[96] && f[545];
	
	// Tree 485, Classifier 5, Iteration: 48
	assign leaf[6939] = !f[264] && !f[241] && !f[239] && !f[243];
	assign leaf[6940] = !f[264] && !f[241] && !f[239] && f[243];
	assign leaf[6941] = !f[264] && !f[241] && f[239] && !f[187];
	assign leaf[6942] = !f[264] && !f[241] && f[239] && f[187];
	assign leaf[6943] = !f[264] && f[241] && !f[217] && !f[238];
	assign leaf[6944] = !f[264] && f[241] && !f[217] && f[238];
	assign leaf[6945] = !f[264] && f[241] && f[217] && !f[239];
	assign leaf[6946] = !f[264] && f[241] && f[217] && f[239];
	assign leaf[6947] = f[264] && !f[241] && !f[157] && !f[296];
	assign leaf[6948] = f[264] && !f[241] && !f[157] && f[296];
	assign leaf[6949] = f[264] && !f[241] && f[157] && !f[244];
	assign leaf[6950] = f[264] && !f[241] && f[157] && f[244];
	assign leaf[6951] = f[264] && f[241] && !f[352] && !f[543];
	assign leaf[6952] = f[264] && f[241] && !f[352] && f[543];
	assign leaf[6953] = f[264] && f[241] && f[352] && !f[243];
	assign leaf[6954] = f[264] && f[241] && f[352] && f[243];
	
	// Tree 486, Classifier 6, Iteration: 48
	assign leaf[6955] = !f[163] && !f[269] && !f[295] && !f[185];
	assign leaf[6956] = !f[163] && !f[269] && !f[295] && f[185];
	assign leaf[6957] = !f[163] && !f[269] && f[295] && !f[185];
	assign leaf[6958] = !f[163] && !f[269] && f[295] && f[185];
	assign leaf[6959] = !f[163] && f[269] && !f[350] && !f[525];
	assign leaf[6960] = !f[163] && f[269] && !f[350] && f[525];
	assign leaf[6961] = !f[163] && f[269] && f[350] && !f[380];
	assign leaf[6962] = !f[163] && f[269] && f[350] && f[380];
	assign leaf[6963] = f[163] && !f[328] && !f[492] && !f[515];
	assign leaf[6964] = f[163] && !f[328] && !f[492] && f[515];
	assign leaf[6965] = f[163] && !f[328] && f[492] && !f[220];
	assign leaf[6966] = f[163] && !f[328] && f[492] && f[220];
	assign leaf[6967] = f[163] && f[328];
	
	// Tree 487, Classifier 7, Iteration: 48
	assign leaf[6968] = !f[128] && !f[296] && !f[431] && !f[485];
	assign leaf[6969] = !f[128] && !f[296] && !f[431] && f[485];
	assign leaf[6970] = !f[128] && !f[296] && f[431] && !f[457];
	assign leaf[6971] = !f[128] && !f[296] && f[431] && f[457];
	assign leaf[6972] = !f[128] && f[296] && !f[404] && !f[492];
	assign leaf[6973] = !f[128] && f[296] && !f[404] && f[492];
	assign leaf[6974] = !f[128] && f[296] && f[404] && !f[318];
	assign leaf[6975] = !f[128] && f[296] && f[404] && f[318];
	assign leaf[6976] = f[128];
	
	// Tree 488, Classifier 8, Iteration: 48
	assign leaf[6977] = !f[273] && !f[289] && !f[375] && !f[320];
	assign leaf[6978] = !f[273] && !f[289] && !f[375] && f[320];
	assign leaf[6979] = !f[273] && !f[289] && f[375] && !f[315];
	assign leaf[6980] = !f[273] && !f[289] && f[375] && f[315];
	assign leaf[6981] = !f[273] && f[289] && !f[375] && !f[320];
	assign leaf[6982] = !f[273] && f[289] && !f[375] && f[320];
	assign leaf[6983] = !f[273] && f[289] && f[375] && !f[401];
	assign leaf[6984] = !f[273] && f[289] && f[375] && f[401];
	assign leaf[6985] = f[273] && !f[322] && !f[402] && !f[348];
	assign leaf[6986] = f[273] && !f[322] && !f[402] && f[348];
	assign leaf[6987] = f[273] && !f[322] && f[402] && !f[288];
	assign leaf[6988] = f[273] && !f[322] && f[402] && f[288];
	assign leaf[6989] = f[273] && f[322] && !f[347] && !f[261];
	assign leaf[6990] = f[273] && f[322] && !f[347] && f[261];
	assign leaf[6991] = f[273] && f[322] && f[347] && !f[519];
	assign leaf[6992] = f[273] && f[322] && f[347] && f[519];
	
	// Tree 489, Classifier 9, Iteration: 48
	assign leaf[6993] = !f[162] && !f[175] && !f[229] && !f[720];
	assign leaf[6994] = !f[162] && !f[175] && !f[229] && f[720];
	assign leaf[6995] = !f[162] && !f[175] && f[229] && !f[369];
	assign leaf[6996] = !f[162] && !f[175] && f[229] && f[369];
	assign leaf[6997] = !f[162] && f[175] && !f[257] && !f[353];
	assign leaf[6998] = !f[162] && f[175] && !f[257] && f[353];
	assign leaf[6999] = !f[162] && f[175] && f[257] && !f[266];
	assign leaf[7000] = !f[162] && f[175] && f[257] && f[266];
	assign leaf[7001] = f[162];
	
	// Tree 490, Classifier 0, Iteration: 49
	assign leaf[7002] = !f[414] && !f[382] && !f[516] && !f[655];
	assign leaf[7003] = !f[414] && !f[382] && !f[516] && f[655];
	assign leaf[7004] = !f[414] && !f[382] && f[516] && !f[151];
	assign leaf[7005] = !f[414] && !f[382] && f[516] && f[151];
	assign leaf[7006] = !f[414] && f[382] && !f[403] && !f[373];
	assign leaf[7007] = !f[414] && f[382] && !f[403] && f[373];
	assign leaf[7008] = !f[414] && f[382] && f[403] && !f[380];
	assign leaf[7009] = !f[414] && f[382] && f[403] && f[380];
	assign leaf[7010] = f[414] && !f[190] && !f[329] && !f[273];
	assign leaf[7011] = f[414] && !f[190] && !f[329] && f[273];
	assign leaf[7012] = f[414] && !f[190] && f[329] && !f[513];
	assign leaf[7013] = f[414] && !f[190] && f[329] && f[513];
	assign leaf[7014] = f[414] && f[190] && !f[521];
	assign leaf[7015] = f[414] && f[190] && f[521] && !f[492];
	assign leaf[7016] = f[414] && f[190] && f[521] && f[492];
	
	// Tree 491, Classifier 1, Iteration: 49
	assign leaf[7017] = !f[556] && !f[260] && !f[552] && !f[99];
	assign leaf[7018] = !f[556] && !f[260] && !f[552] && f[99];
	assign leaf[7019] = !f[556] && !f[260] && f[552] && !f[433];
	assign leaf[7020] = !f[556] && !f[260] && f[552] && f[433];
	assign leaf[7021] = !f[556] && f[260] && !f[625] && !f[543];
	assign leaf[7022] = !f[556] && f[260] && !f[625] && f[543];
	assign leaf[7023] = !f[556] && f[260] && f[625];
	assign leaf[7024] = f[556];
	
	// Tree 492, Classifier 2, Iteration: 49
	assign leaf[7025] = !f[104] && !f[70] && !f[445] && !f[501];
	assign leaf[7026] = !f[104] && !f[70] && !f[445] && f[501];
	assign leaf[7027] = !f[104] && !f[70] && f[445] && !f[552];
	assign leaf[7028] = !f[104] && !f[70] && f[445] && f[552];
	assign leaf[7029] = !f[104] && f[70] && !f[152] && !f[493];
	assign leaf[7030] = !f[104] && f[70] && !f[152] && f[493];
	assign leaf[7031] = !f[104] && f[70] && f[152];
	assign leaf[7032] = f[104] && !f[431] && !f[324];
	assign leaf[7033] = f[104] && !f[431] && f[324];
	assign leaf[7034] = f[104] && f[431] && !f[322];
	assign leaf[7035] = f[104] && f[431] && f[322];
	
	// Tree 493, Classifier 3, Iteration: 49
	assign leaf[7036] = !f[228] && !f[406] && !f[96] && !f[436];
	assign leaf[7037] = !f[228] && !f[406] && !f[96] && f[436];
	assign leaf[7038] = !f[228] && !f[406] && f[96] && !f[431];
	assign leaf[7039] = !f[228] && !f[406] && f[96] && f[431];
	assign leaf[7040] = !f[228] && f[406] && !f[287] && !f[181];
	assign leaf[7041] = !f[228] && f[406] && !f[287] && f[181];
	assign leaf[7042] = !f[228] && f[406] && f[287] && !f[262];
	assign leaf[7043] = !f[228] && f[406] && f[287] && f[262];
	assign leaf[7044] = f[228] && !f[375] && !f[439] && !f[630];
	assign leaf[7045] = f[228] && !f[375] && !f[439] && f[630];
	assign leaf[7046] = f[228] && !f[375] && f[439] && !f[212];
	assign leaf[7047] = f[228] && !f[375] && f[439] && f[212];
	assign leaf[7048] = f[228] && f[375] && !f[344] && !f[293];
	assign leaf[7049] = f[228] && f[375] && !f[344] && f[293];
	assign leaf[7050] = f[228] && f[375] && f[344];
	
	// Tree 494, Classifier 4, Iteration: 49
	assign leaf[7051] = !f[93] && !f[520] && !f[632] && !f[385];
	assign leaf[7052] = !f[93] && !f[520] && !f[632] && f[385];
	assign leaf[7053] = !f[93] && !f[520] && f[632] && !f[485];
	assign leaf[7054] = !f[93] && !f[520] && f[632] && f[485];
	assign leaf[7055] = !f[93] && f[520] && !f[628] && !f[236];
	assign leaf[7056] = !f[93] && f[520] && !f[628] && f[236];
	assign leaf[7057] = !f[93] && f[520] && f[628] && !f[241];
	assign leaf[7058] = !f[93] && f[520] && f[628] && f[241];
	assign leaf[7059] = f[93] && !f[456];
	assign leaf[7060] = f[93] && f[456];
	
	// Tree 495, Classifier 5, Iteration: 49
	assign leaf[7061] = !f[411] && !f[329] && !f[325] && !f[215];
	assign leaf[7062] = !f[411] && !f[329] && !f[325] && f[215];
	assign leaf[7063] = !f[411] && !f[329] && f[325] && !f[352];
	assign leaf[7064] = !f[411] && !f[329] && f[325] && f[352];
	assign leaf[7065] = !f[411] && f[329] && !f[245] && !f[440];
	assign leaf[7066] = !f[411] && f[329] && !f[245] && f[440];
	assign leaf[7067] = !f[411] && f[329] && f[245] && !f[247];
	assign leaf[7068] = !f[411] && f[329] && f[245] && f[247];
	assign leaf[7069] = f[411] && !f[329] && !f[179] && !f[237];
	assign leaf[7070] = f[411] && !f[329] && !f[179] && f[237];
	assign leaf[7071] = f[411] && !f[329] && f[179] && !f[130];
	assign leaf[7072] = f[411] && !f[329] && f[179] && f[130];
	assign leaf[7073] = f[411] && f[329] && !f[150] && !f[130];
	assign leaf[7074] = f[411] && f[329] && !f[150] && f[130];
	assign leaf[7075] = f[411] && f[329] && f[150];
	
	// Tree 496, Classifier 6, Iteration: 49
	assign leaf[7076] = !f[299] && !f[301] && !f[245] && !f[324];
	assign leaf[7077] = !f[299] && !f[301] && !f[245] && f[324];
	assign leaf[7078] = !f[299] && !f[301] && f[245] && !f[541];
	assign leaf[7079] = !f[299] && !f[301] && f[245] && f[541];
	assign leaf[7080] = !f[299] && f[301] && !f[260];
	assign leaf[7081] = !f[299] && f[301] && f[260] && !f[358];
	assign leaf[7082] = !f[299] && f[301] && f[260] && f[358];
	assign leaf[7083] = f[299] && !f[382] && !f[512] && !f[149];
	assign leaf[7084] = f[299] && !f[382] && !f[512] && f[149];
	assign leaf[7085] = f[299] && !f[382] && f[512] && !f[571];
	assign leaf[7086] = f[299] && !f[382] && f[512] && f[571];
	assign leaf[7087] = f[299] && f[382] && !f[357] && !f[456];
	assign leaf[7088] = f[299] && f[382] && !f[357] && f[456];
	assign leaf[7089] = f[299] && f[382] && f[357] && !f[383];
	assign leaf[7090] = f[299] && f[382] && f[357] && f[383];
	
	// Tree 497, Classifier 7, Iteration: 49
	assign leaf[7091] = !f[125] && !f[244] && !f[527] && !f[324];
	assign leaf[7092] = !f[125] && !f[244] && !f[527] && f[324];
	assign leaf[7093] = !f[125] && !f[244] && f[527] && !f[404];
	assign leaf[7094] = !f[125] && !f[244] && f[527] && f[404];
	assign leaf[7095] = !f[125] && f[244] && !f[604] && !f[207];
	assign leaf[7096] = !f[125] && f[244] && !f[604] && f[207];
	assign leaf[7097] = !f[125] && f[244] && f[604] && !f[494];
	assign leaf[7098] = !f[125] && f[244] && f[604] && f[494];
	assign leaf[7099] = f[125] && !f[486];
	assign leaf[7100] = f[125] && f[486];
	
	// Tree 498, Classifier 8, Iteration: 49
	assign leaf[7101] = !f[441] && !f[678] && !f[289] && !f[375];
	assign leaf[7102] = !f[441] && !f[678] && !f[289] && f[375];
	assign leaf[7103] = !f[441] && !f[678] && f[289] && !f[545];
	assign leaf[7104] = !f[441] && !f[678] && f[289] && f[545];
	assign leaf[7105] = !f[441] && f[678] && !f[512] && !f[406];
	assign leaf[7106] = !f[441] && f[678] && !f[512] && f[406];
	assign leaf[7107] = !f[441] && f[678] && f[512] && !f[566];
	assign leaf[7108] = !f[441] && f[678] && f[512] && f[566];
	assign leaf[7109] = f[441] && !f[523] && !f[411] && !f[596];
	assign leaf[7110] = f[441] && !f[523] && !f[411] && f[596];
	assign leaf[7111] = f[441] && !f[523] && f[411] && !f[160];
	assign leaf[7112] = f[441] && !f[523] && f[411] && f[160];
	assign leaf[7113] = f[441] && f[523] && !f[218] && !f[214];
	assign leaf[7114] = f[441] && f[523] && !f[218] && f[214];
	assign leaf[7115] = f[441] && f[523] && f[218] && !f[239];
	assign leaf[7116] = f[441] && f[523] && f[218] && f[239];
	
	// Tree 499, Classifier 9, Iteration: 49
	assign leaf[7117] = !f[573] && !f[711] && !f[404] && !f[461];
	assign leaf[7118] = !f[573] && !f[711] && !f[404] && f[461];
	assign leaf[7119] = !f[573] && !f[711] && f[404] && !f[456];
	assign leaf[7120] = !f[573] && !f[711] && f[404] && f[456];
	assign leaf[7121] = !f[573] && f[711] && !f[412] && !f[600];
	assign leaf[7122] = !f[573] && f[711] && !f[412] && f[600];
	assign leaf[7123] = !f[573] && f[711] && f[412] && !f[494];
	assign leaf[7124] = !f[573] && f[711] && f[412] && f[494];
	assign leaf[7125] = f[573] && !f[207] && !f[549] && !f[489];
	assign leaf[7126] = f[573] && !f[207] && !f[549] && f[489];
	assign leaf[7127] = f[573] && !f[207] && f[549] && !f[484];
	assign leaf[7128] = f[573] && !f[207] && f[549] && f[484];
	assign leaf[7129] = f[573] && f[207] && !f[489] && !f[458];
	assign leaf[7130] = f[573] && f[207] && !f[489] && f[458];
	assign leaf[7131] = f[573] && f[207] && f[489] && !f[290];
	assign leaf[7132] = f[573] && f[207] && f[489] && f[290];
	
	// Tree 500, Classifier 0, Iteration: 50
	assign leaf[7133] = !f[572] && !f[460] && !f[404] && !f[537];
	assign leaf[7134] = !f[572] && !f[460] && !f[404] && f[537];
	assign leaf[7135] = !f[572] && !f[460] && f[404] && !f[266];
	assign leaf[7136] = !f[572] && !f[460] && f[404] && f[266];
	assign leaf[7137] = !f[572] && f[460] && !f[570] && !f[189];
	assign leaf[7138] = !f[572] && f[460] && !f[570] && f[189];
	assign leaf[7139] = !f[572] && f[460] && f[570] && !f[628];
	assign leaf[7140] = !f[572] && f[460] && f[570] && f[628];
	assign leaf[7141] = f[572] && !f[683] && !f[596] && !f[241];
	assign leaf[7142] = f[572] && !f[683] && !f[596] && f[241];
	assign leaf[7143] = f[572] && !f[683] && f[596] && !f[245];
	assign leaf[7144] = f[572] && !f[683] && f[596] && f[245];
	assign leaf[7145] = f[572] && f[683] && !f[577];
	assign leaf[7146] = f[572] && f[683] && f[577];
	
	// Tree 501, Classifier 1, Iteration: 50
	assign leaf[7147] = !f[96] && !f[608] && !f[510] && !f[289];
	assign leaf[7148] = !f[96] && !f[608] && !f[510] && f[289];
	assign leaf[7149] = !f[96] && !f[608] && f[510];
	assign leaf[7150] = !f[96] && f[608] && !f[488] && !f[295];
	assign leaf[7151] = !f[96] && f[608] && !f[488] && f[295];
	assign leaf[7152] = !f[96] && f[608] && f[488] && !f[238];
	assign leaf[7153] = !f[96] && f[608] && f[488] && f[238];
	assign leaf[7154] = f[96] && !f[182];
	assign leaf[7155] = f[96] && f[182];
	
	// Tree 502, Classifier 2, Iteration: 50
	assign leaf[7156] = !f[95] && !f[390] && !f[235] && !f[351];
	assign leaf[7157] = !f[95] && !f[390] && !f[235] && f[351];
	assign leaf[7158] = !f[95] && !f[390] && f[235] && !f[401];
	assign leaf[7159] = !f[95] && !f[390] && f[235] && f[401];
	assign leaf[7160] = !f[95] && f[390];
	assign leaf[7161] = f[95] && !f[262] && !f[453] && !f[402];
	assign leaf[7162] = f[95] && !f[262] && !f[453] && f[402];
	assign leaf[7163] = f[95] && !f[262] && f[453];
	assign leaf[7164] = f[95] && f[262];
	
	// Tree 503, Classifier 3, Iteration: 50
	assign leaf[7165] = !f[429] && !f[544] && !f[489] && !f[459];
	assign leaf[7166] = !f[429] && !f[544] && !f[489] && f[459];
	assign leaf[7167] = !f[429] && !f[544] && f[489] && !f[460];
	assign leaf[7168] = !f[429] && !f[544] && f[489] && f[460];
	assign leaf[7169] = !f[429] && f[544] && !f[538] && !f[572];
	assign leaf[7170] = !f[429] && f[544] && !f[538] && f[572];
	assign leaf[7171] = !f[429] && f[544] && f[538] && !f[294];
	assign leaf[7172] = !f[429] && f[544] && f[538] && f[294];
	assign leaf[7173] = f[429] && !f[460] && !f[484] && !f[405];
	assign leaf[7174] = f[429] && !f[460] && !f[484] && f[405];
	assign leaf[7175] = f[429] && !f[460] && f[484] && !f[402];
	assign leaf[7176] = f[429] && !f[460] && f[484] && f[402];
	assign leaf[7177] = f[429] && f[460] && !f[349] && !f[438];
	assign leaf[7178] = f[429] && f[460] && !f[349] && f[438];
	assign leaf[7179] = f[429] && f[460] && f[349] && !f[657];
	assign leaf[7180] = f[429] && f[460] && f[349] && f[657];
	
	// Tree 504, Classifier 4, Iteration: 50
	assign leaf[7181] = !f[286] && !f[184] && !f[240] && !f[323];
	assign leaf[7182] = !f[286] && !f[184] && !f[240] && f[323];
	assign leaf[7183] = !f[286] && !f[184] && f[240] && !f[238];
	assign leaf[7184] = !f[286] && !f[184] && f[240] && f[238];
	assign leaf[7185] = !f[286] && f[184] && !f[187] && !f[267];
	assign leaf[7186] = !f[286] && f[184] && !f[187] && f[267];
	assign leaf[7187] = !f[286] && f[184] && f[187] && !f[467];
	assign leaf[7188] = !f[286] && f[184] && f[187] && f[467];
	assign leaf[7189] = f[286] && !f[213] && !f[244] && !f[354];
	assign leaf[7190] = f[286] && !f[213] && !f[244] && f[354];
	assign leaf[7191] = f[286] && !f[213] && f[244] && !f[660];
	assign leaf[7192] = f[286] && !f[213] && f[244] && f[660];
	assign leaf[7193] = f[286] && f[213] && !f[205] && !f[687];
	assign leaf[7194] = f[286] && f[213] && !f[205] && f[687];
	assign leaf[7195] = f[286] && f[213] && f[205] && !f[636];
	assign leaf[7196] = f[286] && f[213] && f[205] && f[636];
	
	// Tree 505, Classifier 5, Iteration: 50
	assign leaf[7197] = !f[102] && !f[556] && !f[433] && !f[468];
	assign leaf[7198] = !f[102] && !f[556] && !f[433] && f[468];
	assign leaf[7199] = !f[102] && !f[556] && f[433] && !f[684];
	assign leaf[7200] = !f[102] && !f[556] && f[433] && f[684];
	assign leaf[7201] = !f[102] && f[556] && !f[639] && !f[606];
	assign leaf[7202] = !f[102] && f[556] && !f[639] && f[606];
	assign leaf[7203] = !f[102] && f[556] && f[639];
	assign leaf[7204] = f[102] && !f[604] && !f[404];
	assign leaf[7205] = f[102] && !f[604] && f[404];
	assign leaf[7206] = f[102] && f[604] && !f[344] && !f[349];
	assign leaf[7207] = f[102] && f[604] && !f[344] && f[349];
	assign leaf[7208] = f[102] && f[604] && f[344];
	
	// Tree 506, Classifier 6, Iteration: 50
	assign leaf[7209] = !f[652] && !f[160] && !f[240] && !f[213];
	assign leaf[7210] = !f[652] && !f[160] && !f[240] && f[213];
	assign leaf[7211] = !f[652] && !f[160] && f[240] && !f[158];
	assign leaf[7212] = !f[652] && !f[160] && f[240] && f[158];
	assign leaf[7213] = !f[652] && f[160] && !f[274] && !f[353];
	assign leaf[7214] = !f[652] && f[160] && !f[274] && f[353];
	assign leaf[7215] = !f[652] && f[160] && f[274];
	assign leaf[7216] = f[652] && !f[163];
	assign leaf[7217] = f[652] && f[163];
	
	// Tree 507, Classifier 7, Iteration: 50
	assign leaf[7218] = !f[743] && !f[354] && !f[239] && !f[358];
	assign leaf[7219] = !f[743] && !f[354] && !f[239] && f[358];
	assign leaf[7220] = !f[743] && !f[354] && f[239] && !f[549];
	assign leaf[7221] = !f[743] && !f[354] && f[239] && f[549];
	assign leaf[7222] = !f[743] && f[354] && !f[459] && !f[401];
	assign leaf[7223] = !f[743] && f[354] && !f[459] && f[401];
	assign leaf[7224] = !f[743] && f[354] && f[459] && !f[401];
	assign leaf[7225] = !f[743] && f[354] && f[459] && f[401];
	assign leaf[7226] = f[743] && !f[264] && !f[231] && !f[716];
	assign leaf[7227] = f[743] && !f[264] && !f[231] && f[716];
	assign leaf[7228] = f[743] && !f[264] && f[231];
	assign leaf[7229] = f[743] && f[264] && !f[343] && !f[235];
	assign leaf[7230] = f[743] && f[264] && !f[343] && f[235];
	assign leaf[7231] = f[743] && f[264] && f[343] && !f[260];
	assign leaf[7232] = f[743] && f[264] && f[343] && f[260];
	
	// Tree 508, Classifier 8, Iteration: 50
	assign leaf[7233] = !f[705] && !f[219] && !f[708] && !f[120];
	assign leaf[7234] = !f[705] && !f[219] && !f[708] && f[120];
	assign leaf[7235] = !f[705] && !f[219] && f[708] && !f[568];
	assign leaf[7236] = !f[705] && !f[219] && f[708] && f[568];
	assign leaf[7237] = !f[705] && f[219] && !f[379] && !f[543];
	assign leaf[7238] = !f[705] && f[219] && !f[379] && f[543];
	assign leaf[7239] = !f[705] && f[219] && f[379] && !f[346];
	assign leaf[7240] = !f[705] && f[219] && f[379] && f[346];
	assign leaf[7241] = f[705];
	
	// Tree 509, Classifier 9, Iteration: 50
	assign leaf[7242] = !f[129] && !f[415] && !f[244] && !f[326];
	assign leaf[7243] = !f[129] && !f[415] && !f[244] && f[326];
	assign leaf[7244] = !f[129] && !f[415] && f[244] && !f[330];
	assign leaf[7245] = !f[129] && !f[415] && f[244] && f[330];
	assign leaf[7246] = !f[129] && f[415] && !f[302] && !f[430];
	assign leaf[7247] = !f[129] && f[415] && !f[302] && f[430];
	assign leaf[7248] = !f[129] && f[415] && f[302] && !f[403];
	assign leaf[7249] = !f[129] && f[415] && f[302] && f[403];
	assign leaf[7250] = f[129] && !f[217] && !f[185];
	assign leaf[7251] = f[129] && !f[217] && f[185];
	assign leaf[7252] = f[129] && f[217];
	
	// Tree 510, Classifier 0, Iteration: 51
	assign leaf[7253] = !f[133] && !f[397] && !f[428] && !f[567];
	assign leaf[7254] = !f[133] && !f[397] && !f[428] && f[567];
	assign leaf[7255] = !f[133] && !f[397] && f[428] && !f[458];
	assign leaf[7256] = !f[133] && !f[397] && f[428] && f[458];
	assign leaf[7257] = !f[133] && f[397] && !f[626] && !f[498];
	assign leaf[7258] = !f[133] && f[397] && !f[626] && f[498];
	assign leaf[7259] = !f[133] && f[397] && f[626] && !f[430];
	assign leaf[7260] = !f[133] && f[397] && f[626] && f[430];
	assign leaf[7261] = f[133] && !f[653] && !f[516];
	assign leaf[7262] = f[133] && !f[653] && f[516];
	assign leaf[7263] = f[133] && f[653] && !f[512];
	assign leaf[7264] = f[133] && f[653] && f[512];
	
	// Tree 511, Classifier 1, Iteration: 51
	assign leaf[7265] = !f[604] && !f[180] && !f[264] && !f[296];
	assign leaf[7266] = !f[604] && !f[180] && !f[264] && f[296];
	assign leaf[7267] = !f[604] && !f[180] && f[264] && !f[663];
	assign leaf[7268] = !f[604] && !f[180] && f[264] && f[663];
	assign leaf[7269] = !f[604] && f[180] && !f[269] && !f[125];
	assign leaf[7270] = !f[604] && f[180] && !f[269] && f[125];
	assign leaf[7271] = !f[604] && f[180] && f[269] && !f[152];
	assign leaf[7272] = !f[604] && f[180] && f[269] && f[152];
	assign leaf[7273] = f[604] && !f[546] && !f[460] && !f[658];
	assign leaf[7274] = f[604] && !f[546] && !f[460] && f[658];
	assign leaf[7275] = f[604] && !f[546] && f[460] && !f[576];
	assign leaf[7276] = f[604] && !f[546] && f[460] && f[576];
	assign leaf[7277] = f[604] && f[546] && !f[514] && !f[595];
	assign leaf[7278] = f[604] && f[546] && !f[514] && f[595];
	assign leaf[7279] = f[604] && f[546] && f[514] && !f[291];
	assign leaf[7280] = f[604] && f[546] && f[514] && f[291];
	
	// Tree 512, Classifier 2, Iteration: 51
	assign leaf[7281] = !f[134] && !f[411] && !f[356] && !f[470];
	assign leaf[7282] = !f[134] && !f[411] && !f[356] && f[470];
	assign leaf[7283] = !f[134] && !f[411] && f[356] && !f[324];
	assign leaf[7284] = !f[134] && !f[411] && f[356] && f[324];
	assign leaf[7285] = !f[134] && f[411] && !f[493] && !f[524];
	assign leaf[7286] = !f[134] && f[411] && !f[493] && f[524];
	assign leaf[7287] = !f[134] && f[411] && f[493] && !f[515];
	assign leaf[7288] = !f[134] && f[411] && f[493] && f[515];
	assign leaf[7289] = f[134] && !f[301];
	assign leaf[7290] = f[134] && f[301] && !f[467];
	assign leaf[7291] = f[134] && f[301] && f[467];
	
	// Tree 513, Classifier 3, Iteration: 51
	assign leaf[7292] = !f[373] && !f[316] && !f[718] && !f[689];
	assign leaf[7293] = !f[373] && !f[316] && !f[718] && f[689];
	assign leaf[7294] = !f[373] && !f[316] && f[718] && !f[460];
	assign leaf[7295] = !f[373] && !f[316] && f[718] && f[460];
	assign leaf[7296] = !f[373] && f[316] && !f[264] && !f[407];
	assign leaf[7297] = !f[373] && f[316] && !f[264] && f[407];
	assign leaf[7298] = !f[373] && f[316] && f[264] && !f[398];
	assign leaf[7299] = !f[373] && f[316] && f[264] && f[398];
	assign leaf[7300] = f[373] && !f[289] && !f[315] && !f[607];
	assign leaf[7301] = f[373] && !f[289] && !f[315] && f[607];
	assign leaf[7302] = f[373] && !f[289] && f[315] && !f[287];
	assign leaf[7303] = f[373] && !f[289] && f[315] && f[287];
	assign leaf[7304] = f[373] && f[289] && !f[264] && !f[317];
	assign leaf[7305] = f[373] && f[289] && !f[264] && f[317];
	assign leaf[7306] = f[373] && f[289] && f[264] && !f[183];
	assign leaf[7307] = f[373] && f[289] && f[264] && f[183];
	
	// Tree 514, Classifier 4, Iteration: 51
	assign leaf[7308] = !f[397] && !f[346] && !f[348] && !f[344];
	assign leaf[7309] = !f[397] && !f[346] && !f[348] && f[344];
	assign leaf[7310] = !f[397] && !f[346] && f[348] && !f[490];
	assign leaf[7311] = !f[397] && !f[346] && f[348] && f[490];
	assign leaf[7312] = !f[397] && f[346] && !f[400] && !f[212];
	assign leaf[7313] = !f[397] && f[346] && !f[400] && f[212];
	assign leaf[7314] = !f[397] && f[346] && f[400] && !f[243];
	assign leaf[7315] = !f[397] && f[346] && f[400] && f[243];
	assign leaf[7316] = f[397] && !f[359] && !f[379] && !f[323];
	assign leaf[7317] = f[397] && !f[359] && !f[379] && f[323];
	assign leaf[7318] = f[397] && !f[359] && f[379] && !f[372];
	assign leaf[7319] = f[397] && !f[359] && f[379] && f[372];
	assign leaf[7320] = f[397] && f[359] && !f[429];
	assign leaf[7321] = f[397] && f[359] && f[429];
	
	// Tree 515, Classifier 5, Iteration: 51
	assign leaf[7322] = !f[200] && !f[717] && !f[599] && !f[681];
	assign leaf[7323] = !f[200] && !f[717] && !f[599] && f[681];
	assign leaf[7324] = !f[200] && !f[717] && f[599] && !f[602];
	assign leaf[7325] = !f[200] && !f[717] && f[599] && f[602];
	assign leaf[7326] = !f[200] && f[717] && !f[577] && !f[657];
	assign leaf[7327] = !f[200] && f[717] && !f[577] && f[657];
	assign leaf[7328] = !f[200] && f[717] && f[577] && !f[214];
	assign leaf[7329] = !f[200] && f[717] && f[577] && f[214];
	assign leaf[7330] = f[200];
	
	// Tree 516, Classifier 6, Iteration: 51
	assign leaf[7331] = !f[428] && !f[235] && !f[124] && !f[567];
	assign leaf[7332] = !f[428] && !f[235] && !f[124] && f[567];
	assign leaf[7333] = !f[428] && !f[235] && f[124] && !f[426];
	assign leaf[7334] = !f[428] && !f[235] && f[124] && f[426];
	assign leaf[7335] = !f[428] && f[235] && !f[96] && !f[98];
	assign leaf[7336] = !f[428] && f[235] && !f[96] && f[98];
	assign leaf[7337] = !f[428] && f[235] && f[96] && !f[599];
	assign leaf[7338] = !f[428] && f[235] && f[96] && f[599];
	assign leaf[7339] = f[428] && !f[541] && !f[236] && !f[548];
	assign leaf[7340] = f[428] && !f[541] && !f[236] && f[548];
	assign leaf[7341] = f[428] && !f[541] && f[236] && !f[151];
	assign leaf[7342] = f[428] && !f[541] && f[236] && f[151];
	assign leaf[7343] = f[428] && f[541] && !f[318] && !f[264];
	assign leaf[7344] = f[428] && f[541] && !f[318] && f[264];
	assign leaf[7345] = f[428] && f[541] && f[318] && !f[157];
	assign leaf[7346] = f[428] && f[541] && f[318] && f[157];
	
	// Tree 517, Classifier 7, Iteration: 51
	assign leaf[7347] = !f[690] && !f[634] && !f[177] && !f[232];
	assign leaf[7348] = !f[690] && !f[634] && !f[177] && f[232];
	assign leaf[7349] = !f[690] && !f[634] && f[177] && !f[523];
	assign leaf[7350] = !f[690] && !f[634] && f[177] && f[523];
	assign leaf[7351] = !f[690] && f[634] && !f[434] && !f[342];
	assign leaf[7352] = !f[690] && f[634] && !f[434] && f[342];
	assign leaf[7353] = !f[690] && f[634] && f[434] && !f[468];
	assign leaf[7354] = !f[690] && f[634] && f[434] && f[468];
	assign leaf[7355] = f[690] && !f[291] && !f[522] && !f[633];
	assign leaf[7356] = f[690] && !f[291] && !f[522] && f[633];
	assign leaf[7357] = f[690] && !f[291] && f[522] && !f[496];
	assign leaf[7358] = f[690] && !f[291] && f[522] && f[496];
	assign leaf[7359] = f[690] && f[291] && !f[489] && !f[686];
	assign leaf[7360] = f[690] && f[291] && !f[489] && f[686];
	assign leaf[7361] = f[690] && f[291] && f[489] && !f[286];
	assign leaf[7362] = f[690] && f[291] && f[489] && f[286];
	
	// Tree 518, Classifier 8, Iteration: 51
	assign leaf[7363] = !f[452] && !f[333] && !f[705] && !f[563];
	assign leaf[7364] = !f[452] && !f[333] && !f[705] && f[563];
	assign leaf[7365] = !f[452] && !f[333] && f[705];
	assign leaf[7366] = !f[452] && f[333] && !f[299] && !f[573];
	assign leaf[7367] = !f[452] && f[333] && !f[299] && f[573];
	assign leaf[7368] = !f[452] && f[333] && f[299];
	assign leaf[7369] = f[452];
	
	// Tree 519, Classifier 9, Iteration: 51
	assign leaf[7370] = !f[340] && !f[353] && !f[385] && !f[156];
	assign leaf[7371] = !f[340] && !f[353] && !f[385] && f[156];
	assign leaf[7372] = !f[340] && !f[353] && f[385] && !f[214];
	assign leaf[7373] = !f[340] && !f[353] && f[385] && f[214];
	assign leaf[7374] = !f[340] && f[353] && !f[574] && !f[712];
	assign leaf[7375] = !f[340] && f[353] && !f[574] && f[712];
	assign leaf[7376] = !f[340] && f[353] && f[574] && !f[543];
	assign leaf[7377] = !f[340] && f[353] && f[574] && f[543];
	assign leaf[7378] = f[340] && !f[346] && !f[688] && !f[526];
	assign leaf[7379] = f[340] && !f[346] && !f[688] && f[526];
	assign leaf[7380] = f[340] && !f[346] && f[688];
	assign leaf[7381] = f[340] && f[346] && !f[214];
	assign leaf[7382] = f[340] && f[346] && f[214];
	
	// Tree 520, Classifier 0, Iteration: 52
	assign leaf[7383] = !f[378] && !f[352] && !f[453] && !f[518];
	assign leaf[7384] = !f[378] && !f[352] && !f[453] && f[518];
	assign leaf[7385] = !f[378] && !f[352] && f[453] && !f[661];
	assign leaf[7386] = !f[378] && !f[352] && f[453] && f[661];
	assign leaf[7387] = !f[378] && f[352] && !f[431] && !f[320];
	assign leaf[7388] = !f[378] && f[352] && !f[431] && f[320];
	assign leaf[7389] = !f[378] && f[352] && f[431] && !f[294];
	assign leaf[7390] = !f[378] && f[352] && f[431] && f[294];
	assign leaf[7391] = f[378] && !f[488] && !f[352] && !f[329];
	assign leaf[7392] = f[378] && !f[488] && !f[352] && f[329];
	assign leaf[7393] = f[378] && !f[488] && f[352] && !f[377];
	assign leaf[7394] = f[378] && !f[488] && f[352] && f[377];
	assign leaf[7395] = f[378] && f[488] && !f[686] && !f[542];
	assign leaf[7396] = f[378] && f[488] && !f[686] && f[542];
	assign leaf[7397] = f[378] && f[488] && f[686];
	
	// Tree 521, Classifier 1, Iteration: 52
	assign leaf[7398] = !f[72] && !f[493] && !f[148] && !f[244];
	assign leaf[7399] = !f[72] && !f[493] && !f[148] && f[244];
	assign leaf[7400] = !f[72] && !f[493] && f[148] && !f[570];
	assign leaf[7401] = !f[72] && !f[493] && f[148] && f[570];
	assign leaf[7402] = !f[72] && f[493] && !f[576] && !f[179];
	assign leaf[7403] = !f[72] && f[493] && !f[576] && f[179];
	assign leaf[7404] = !f[72] && f[493] && f[576] && !f[519];
	assign leaf[7405] = !f[72] && f[493] && f[576] && f[519];
	assign leaf[7406] = f[72];
	
	// Tree 522, Classifier 2, Iteration: 52
	assign leaf[7407] = !f[708] && !f[514] && !f[432] && !f[231];
	assign leaf[7408] = !f[708] && !f[514] && !f[432] && f[231];
	assign leaf[7409] = !f[708] && !f[514] && f[432] && !f[408];
	assign leaf[7410] = !f[708] && !f[514] && f[432] && f[408];
	assign leaf[7411] = !f[708] && f[514] && !f[597] && !f[287];
	assign leaf[7412] = !f[708] && f[514] && !f[597] && f[287];
	assign leaf[7413] = !f[708] && f[514] && f[597] && !f[184];
	assign leaf[7414] = !f[708] && f[514] && f[597] && f[184];
	assign leaf[7415] = f[708] && !f[460];
	assign leaf[7416] = f[708] && f[460];
	
	// Tree 523, Classifier 3, Iteration: 52
	assign leaf[7417] = !f[401] && !f[716] && !f[459] && !f[537];
	assign leaf[7418] = !f[401] && !f[716] && !f[459] && f[537];
	assign leaf[7419] = !f[401] && !f[716] && f[459] && !f[570];
	assign leaf[7420] = !f[401] && !f[716] && f[459] && f[570];
	assign leaf[7421] = !f[401] && f[716] && !f[433] && !f[576];
	assign leaf[7422] = !f[401] && f[716] && !f[433] && f[576];
	assign leaf[7423] = !f[401] && f[716] && f[433] && !f[347];
	assign leaf[7424] = !f[401] && f[716] && f[433] && f[347];
	assign leaf[7425] = f[401] && !f[482] && !f[344] && !f[513];
	assign leaf[7426] = f[401] && !f[482] && !f[344] && f[513];
	assign leaf[7427] = f[401] && !f[482] && f[344] && !f[347];
	assign leaf[7428] = f[401] && !f[482] && f[344] && f[347];
	assign leaf[7429] = f[401] && f[482] && !f[538] && !f[578];
	assign leaf[7430] = f[401] && f[482] && !f[538] && f[578];
	assign leaf[7431] = f[401] && f[482] && f[538] && !f[541];
	assign leaf[7432] = f[401] && f[482] && f[538] && f[541];
	
	// Tree 524, Classifier 4, Iteration: 52
	assign leaf[7433] = !f[347] && !f[344] && !f[405] && !f[349];
	assign leaf[7434] = !f[347] && !f[344] && !f[405] && f[349];
	assign leaf[7435] = !f[347] && !f[344] && f[405] && !f[318];
	assign leaf[7436] = !f[347] && !f[344] && f[405] && f[318];
	assign leaf[7437] = !f[347] && f[344] && !f[180] && !f[264];
	assign leaf[7438] = !f[347] && f[344] && !f[180] && f[264];
	assign leaf[7439] = !f[347] && f[344] && f[180] && !f[661];
	assign leaf[7440] = !f[347] && f[344] && f[180] && f[661];
	assign leaf[7441] = f[347] && !f[341] && !f[542] && !f[240];
	assign leaf[7442] = f[347] && !f[341] && !f[542] && f[240];
	assign leaf[7443] = f[347] && !f[341] && f[542] && !f[526];
	assign leaf[7444] = f[347] && !f[341] && f[542] && f[526];
	assign leaf[7445] = f[347] && f[341] && !f[636] && !f[271];
	assign leaf[7446] = f[347] && f[341] && !f[636] && f[271];
	assign leaf[7447] = f[347] && f[341] && f[636];
	
	// Tree 525, Classifier 5, Iteration: 52
	assign leaf[7448] = !f[264] && !f[241] && !f[243] && !f[239];
	assign leaf[7449] = !f[264] && !f[241] && !f[243] && f[239];
	assign leaf[7450] = !f[264] && !f[241] && f[243] && !f[268];
	assign leaf[7451] = !f[264] && !f[241] && f[243] && f[268];
	assign leaf[7452] = !f[264] && f[241] && !f[155] && !f[158];
	assign leaf[7453] = !f[264] && f[241] && !f[155] && f[158];
	assign leaf[7454] = !f[264] && f[241] && f[155] && !f[238];
	assign leaf[7455] = !f[264] && f[241] && f[155] && f[238];
	assign leaf[7456] = f[264] && !f[207] && !f[321] && !f[184];
	assign leaf[7457] = f[264] && !f[207] && !f[321] && f[184];
	assign leaf[7458] = f[264] && !f[207] && f[321] && !f[633];
	assign leaf[7459] = f[264] && !f[207] && f[321] && f[633];
	assign leaf[7460] = f[264] && f[207] && !f[174] && !f[358];
	assign leaf[7461] = f[264] && f[207] && !f[174] && f[358];
	assign leaf[7462] = f[264] && f[207] && f[174] && !f[413];
	assign leaf[7463] = f[264] && f[207] && f[174] && f[413];
	
	// Tree 526, Classifier 6, Iteration: 52
	assign leaf[7464] = !f[409] && !f[98] && !f[571] && !f[323];
	assign leaf[7465] = !f[409] && !f[98] && !f[571] && f[323];
	assign leaf[7466] = !f[409] && !f[98] && f[571] && !f[271];
	assign leaf[7467] = !f[409] && !f[98] && f[571] && f[271];
	assign leaf[7468] = !f[409] && f[98] && !f[579] && !f[353];
	assign leaf[7469] = !f[409] && f[98] && !f[579] && f[353];
	assign leaf[7470] = !f[409] && f[98] && f[579] && !f[601];
	assign leaf[7471] = !f[409] && f[98] && f[579] && f[601];
	assign leaf[7472] = f[409] && !f[441] && !f[327] && !f[325];
	assign leaf[7473] = f[409] && !f[441] && !f[327] && f[325];
	assign leaf[7474] = f[409] && !f[441] && f[327] && !f[149];
	assign leaf[7475] = f[409] && !f[441] && f[327] && f[149];
	assign leaf[7476] = f[409] && f[441] && !f[377] && !f[270];
	assign leaf[7477] = f[409] && f[441] && !f[377] && f[270];
	assign leaf[7478] = f[409] && f[441] && f[377] && !f[484];
	assign leaf[7479] = f[409] && f[441] && f[377] && f[484];
	
	// Tree 527, Classifier 7, Iteration: 52
	assign leaf[7480] = !f[242] && !f[457] && !f[397] && !f[347];
	assign leaf[7481] = !f[242] && !f[457] && !f[397] && f[347];
	assign leaf[7482] = !f[242] && !f[457] && f[397] && !f[513];
	assign leaf[7483] = !f[242] && !f[457] && f[397] && f[513];
	assign leaf[7484] = !f[242] && f[457] && !f[399] && !f[322];
	assign leaf[7485] = !f[242] && f[457] && !f[399] && f[322];
	assign leaf[7486] = !f[242] && f[457] && f[399] && !f[347];
	assign leaf[7487] = !f[242] && f[457] && f[399] && f[347];
	assign leaf[7488] = f[242] && !f[604] && !f[320] && !f[317];
	assign leaf[7489] = f[242] && !f[604] && !f[320] && f[317];
	assign leaf[7490] = f[242] && !f[604] && f[320] && !f[373];
	assign leaf[7491] = f[242] && !f[604] && f[320] && f[373];
	assign leaf[7492] = f[242] && f[604] && !f[716] && !f[655];
	assign leaf[7493] = f[242] && f[604] && !f[716] && f[655];
	assign leaf[7494] = f[242] && f[604] && f[716] && !f[515];
	assign leaf[7495] = f[242] && f[604] && f[716] && f[515];
	
	// Tree 528, Classifier 8, Iteration: 52
	assign leaf[7496] = !f[304] && !f[708] && !f[322] && !f[462];
	assign leaf[7497] = !f[304] && !f[708] && !f[322] && f[462];
	assign leaf[7498] = !f[304] && !f[708] && f[322] && !f[546];
	assign leaf[7499] = !f[304] && !f[708] && f[322] && f[546];
	assign leaf[7500] = !f[304] && f[708] && !f[568] && !f[630];
	assign leaf[7501] = !f[304] && f[708] && !f[568] && f[630];
	assign leaf[7502] = !f[304] && f[708] && f[568];
	assign leaf[7503] = f[304] && !f[322] && !f[486] && !f[653];
	assign leaf[7504] = f[304] && !f[322] && !f[486] && f[653];
	assign leaf[7505] = f[304] && !f[322] && f[486];
	assign leaf[7506] = f[304] && f[322] && !f[212] && !f[268];
	assign leaf[7507] = f[304] && f[322] && !f[212] && f[268];
	assign leaf[7508] = f[304] && f[322] && f[212] && !f[262];
	assign leaf[7509] = f[304] && f[322] && f[212] && f[262];
	
	// Tree 529, Classifier 9, Iteration: 52
	assign leaf[7510] = !f[584] && !f[500] && !f[740] && !f[326];
	assign leaf[7511] = !f[584] && !f[500] && !f[740] && f[326];
	assign leaf[7512] = !f[584] && !f[500] && f[740] && !f[714];
	assign leaf[7513] = !f[584] && !f[500] && f[740] && f[714];
	assign leaf[7514] = !f[584] && f[500];
	assign leaf[7515] = f[584] && !f[297];
	assign leaf[7516] = f[584] && f[297];
	
	// Tree 530, Classifier 0, Iteration: 53
	assign leaf[7517] = !f[713] && !f[605] && !f[406] && !f[637];
	assign leaf[7518] = !f[713] && !f[605] && !f[406] && f[637];
	assign leaf[7519] = !f[713] && !f[605] && f[406] && !f[216];
	assign leaf[7520] = !f[713] && !f[605] && f[406] && f[216];
	assign leaf[7521] = !f[713] && f[605] && !f[207] && !f[683];
	assign leaf[7522] = !f[713] && f[605] && !f[207] && f[683];
	assign leaf[7523] = !f[713] && f[605] && f[207] && !f[624];
	assign leaf[7524] = !f[713] && f[605] && f[207] && f[624];
	assign leaf[7525] = f[713] && !f[295];
	assign leaf[7526] = f[713] && f[295];
	
	// Tree 531, Classifier 1, Iteration: 53
	assign leaf[7527] = !f[316] && !f[627] && !f[240] && !f[185];
	assign leaf[7528] = !f[316] && !f[627] && !f[240] && f[185];
	assign leaf[7529] = !f[316] && !f[627] && f[240] && !f[151];
	assign leaf[7530] = !f[316] && !f[627] && f[240] && f[151];
	assign leaf[7531] = !f[316] && f[627] && !f[296] && !f[606];
	assign leaf[7532] = !f[316] && f[627] && !f[296] && f[606];
	assign leaf[7533] = !f[316] && f[627] && f[296] && !f[352];
	assign leaf[7534] = !f[316] && f[627] && f[296] && f[352];
	assign leaf[7535] = f[316] && !f[597];
	assign leaf[7536] = f[316] && f[597];
	
	// Tree 532, Classifier 2, Iteration: 53
	assign leaf[7537] = !f[242] && !f[154] && !f[213] && !f[299];
	assign leaf[7538] = !f[242] && !f[154] && !f[213] && f[299];
	assign leaf[7539] = !f[242] && !f[154] && f[213] && !f[355];
	assign leaf[7540] = !f[242] && !f[154] && f[213] && f[355];
	assign leaf[7541] = !f[242] && f[154] && !f[159] && !f[240];
	assign leaf[7542] = !f[242] && f[154] && !f[159] && f[240];
	assign leaf[7543] = !f[242] && f[154] && f[159] && !f[358];
	assign leaf[7544] = !f[242] && f[154] && f[159] && f[358];
	assign leaf[7545] = f[242] && !f[156] && !f[509] && !f[688];
	assign leaf[7546] = f[242] && !f[156] && !f[509] && f[688];
	assign leaf[7547] = f[242] && !f[156] && f[509] && !f[464];
	assign leaf[7548] = f[242] && !f[156] && f[509] && f[464];
	assign leaf[7549] = f[242] && f[156] && !f[597] && !f[408];
	assign leaf[7550] = f[242] && f[156] && !f[597] && f[408];
	assign leaf[7551] = f[242] && f[156] && f[597] && !f[594];
	assign leaf[7552] = f[242] && f[156] && f[597] && f[594];
	
	// Tree 533, Classifier 3, Iteration: 53
	assign leaf[7553] = !f[708] && !f[386] && !f[269] && !f[239];
	assign leaf[7554] = !f[708] && !f[386] && !f[269] && f[239];
	assign leaf[7555] = !f[708] && !f[386] && f[269] && !f[101];
	assign leaf[7556] = !f[708] && !f[386] && f[269] && f[101];
	assign leaf[7557] = !f[708] && f[386] && !f[355];
	assign leaf[7558] = !f[708] && f[386] && f[355] && !f[259];
	assign leaf[7559] = !f[708] && f[386] && f[355] && f[259];
	assign leaf[7560] = f[708] && !f[599] && !f[274] && !f[488];
	assign leaf[7561] = f[708] && !f[599] && !f[274] && f[488];
	assign leaf[7562] = f[708] && !f[599] && f[274];
	assign leaf[7563] = f[708] && f[599] && !f[602];
	assign leaf[7564] = f[708] && f[599] && f[602];
	
	// Tree 534, Classifier 4, Iteration: 53
	assign leaf[7565] = !f[122] && !f[128] && !f[376] && !f[399];
	assign leaf[7566] = !f[122] && !f[128] && !f[376] && f[399];
	assign leaf[7567] = !f[122] && !f[128] && f[376] && !f[408];
	assign leaf[7568] = !f[122] && !f[128] && f[376] && f[408];
	assign leaf[7569] = !f[122] && f[128] && !f[405] && !f[598];
	assign leaf[7570] = !f[122] && f[128] && !f[405] && f[598];
	assign leaf[7571] = !f[122] && f[128] && f[405] && !f[267];
	assign leaf[7572] = !f[122] && f[128] && f[405] && f[267];
	assign leaf[7573] = f[122] && !f[546] && !f[630];
	assign leaf[7574] = f[122] && !f[546] && f[630];
	assign leaf[7575] = f[122] && f[546] && !f[513];
	assign leaf[7576] = f[122] && f[546] && f[513];
	
	// Tree 535, Classifier 5, Iteration: 53
	assign leaf[7577] = !f[228] && !f[101] && !f[565] && !f[481];
	assign leaf[7578] = !f[228] && !f[101] && !f[565] && f[481];
	assign leaf[7579] = !f[228] && !f[101] && f[565] && !f[427];
	assign leaf[7580] = !f[228] && !f[101] && f[565] && f[427];
	assign leaf[7581] = !f[228] && f[101] && !f[242] && !f[441];
	assign leaf[7582] = !f[228] && f[101] && !f[242] && f[441];
	assign leaf[7583] = !f[228] && f[101] && f[242];
	assign leaf[7584] = f[228];
	
	// Tree 536, Classifier 6, Iteration: 53
	assign leaf[7585] = !f[91] && !f[202] && !f[439] && !f[409];
	assign leaf[7586] = !f[91] && !f[202] && !f[439] && f[409];
	assign leaf[7587] = !f[91] && !f[202] && f[439] && !f[403];
	assign leaf[7588] = !f[91] && !f[202] && f[439] && f[403];
	assign leaf[7589] = !f[91] && f[202] && !f[426];
	assign leaf[7590] = !f[91] && f[202] && f[426];
	assign leaf[7591] = f[91];
	
	// Tree 537, Classifier 7, Iteration: 53
	assign leaf[7592] = !f[160] && !f[639] && !f[528] && !f[434];
	assign leaf[7593] = !f[160] && !f[639] && !f[528] && f[434];
	assign leaf[7594] = !f[160] && !f[639] && f[528] && !f[381];
	assign leaf[7595] = !f[160] && !f[639] && f[528] && f[381];
	assign leaf[7596] = !f[160] && f[639];
	assign leaf[7597] = f[160] && !f[182];
	assign leaf[7598] = f[160] && f[182];
	
	// Tree 538, Classifier 8, Iteration: 53
	assign leaf[7599] = !f[649] && !f[708] && !f[434] && !f[429];
	assign leaf[7600] = !f[649] && !f[708] && !f[434] && f[429];
	assign leaf[7601] = !f[649] && !f[708] && f[434] && !f[100];
	assign leaf[7602] = !f[649] && !f[708] && f[434] && f[100];
	assign leaf[7603] = !f[649] && f[708] && !f[513] && !f[575];
	assign leaf[7604] = !f[649] && f[708] && !f[513] && f[575];
	assign leaf[7605] = !f[649] && f[708] && f[513];
	assign leaf[7606] = f[649] && !f[539] && !f[247];
	assign leaf[7607] = f[649] && !f[539] && f[247];
	assign leaf[7608] = f[649] && f[539] && !f[347] && !f[349];
	assign leaf[7609] = f[649] && f[539] && !f[347] && f[349];
	assign leaf[7610] = f[649] && f[539] && f[347];
	
	// Tree 539, Classifier 9, Iteration: 53
	assign leaf[7611] = !f[605] && !f[566] && !f[717] && !f[378];
	assign leaf[7612] = !f[605] && !f[566] && !f[717] && f[378];
	assign leaf[7613] = !f[605] && !f[566] && f[717] && !f[233];
	assign leaf[7614] = !f[605] && !f[566] && f[717] && f[233];
	assign leaf[7615] = !f[605] && f[566] && !f[631];
	assign leaf[7616] = !f[605] && f[566] && f[631];
	assign leaf[7617] = f[605] && !f[546] && !f[180] && !f[236];
	assign leaf[7618] = f[605] && !f[546] && !f[180] && f[236];
	assign leaf[7619] = f[605] && !f[546] && f[180] && !f[265];
	assign leaf[7620] = f[605] && !f[546] && f[180] && f[265];
	assign leaf[7621] = f[605] && f[546] && !f[494] && !f[512];
	assign leaf[7622] = f[605] && f[546] && !f[494] && f[512];
	assign leaf[7623] = f[605] && f[546] && f[494] && !f[469];
	assign leaf[7624] = f[605] && f[546] && f[494] && f[469];
	
	// Tree 540, Classifier 0, Iteration: 54
	assign leaf[7625] = !f[713] && !f[710] && !f[427] && !f[344];
	assign leaf[7626] = !f[713] && !f[710] && !f[427] && f[344];
	assign leaf[7627] = !f[713] && !f[710] && f[427] && !f[345];
	assign leaf[7628] = !f[713] && !f[710] && f[427] && f[345];
	assign leaf[7629] = !f[713] && f[710];
	assign leaf[7630] = f[713] && !f[376];
	assign leaf[7631] = f[713] && f[376];
	
	// Tree 541, Classifier 1, Iteration: 54
	assign leaf[7632] = !f[511] && !f[72] && !f[711] && !f[678];
	assign leaf[7633] = !f[511] && !f[72] && !f[711] && f[678];
	assign leaf[7634] = !f[511] && !f[72] && f[711];
	assign leaf[7635] = !f[511] && f[72];
	assign leaf[7636] = f[511] && !f[430] && !f[349];
	assign leaf[7637] = f[511] && !f[430] && f[349];
	assign leaf[7638] = f[511] && f[430] && !f[186];
	assign leaf[7639] = f[511] && f[430] && f[186];
	
	// Tree 542, Classifier 2, Iteration: 54
	assign leaf[7640] = !f[400] && !f[344] && !f[233] && !f[607];
	assign leaf[7641] = !f[400] && !f[344] && !f[233] && f[607];
	assign leaf[7642] = !f[400] && !f[344] && f[233] && !f[466];
	assign leaf[7643] = !f[400] && !f[344] && f[233] && f[466];
	assign leaf[7644] = !f[400] && f[344] && !f[401] && !f[454];
	assign leaf[7645] = !f[400] && f[344] && !f[401] && f[454];
	assign leaf[7646] = !f[400] && f[344] && f[401] && !f[343];
	assign leaf[7647] = !f[400] && f[344] && f[401] && f[343];
	assign leaf[7648] = f[400] && !f[376] && !f[372] && !f[432];
	assign leaf[7649] = f[400] && !f[376] && !f[372] && f[432];
	assign leaf[7650] = f[400] && !f[376] && f[372] && !f[623];
	assign leaf[7651] = f[400] && !f[376] && f[372] && f[623];
	assign leaf[7652] = f[400] && f[376] && !f[659] && !f[295];
	assign leaf[7653] = f[400] && f[376] && !f[659] && f[295];
	assign leaf[7654] = f[400] && f[376] && f[659] && !f[547];
	assign leaf[7655] = f[400] && f[376] && f[659] && f[547];
	
	// Tree 543, Classifier 3, Iteration: 54
	assign leaf[7656] = !f[712] && !f[370] && !f[480] && !f[678];
	assign leaf[7657] = !f[712] && !f[370] && !f[480] && f[678];
	assign leaf[7658] = !f[712] && !f[370] && f[480] && !f[545];
	assign leaf[7659] = !f[712] && !f[370] && f[480] && f[545];
	assign leaf[7660] = !f[712] && f[370] && !f[286] && !f[492];
	assign leaf[7661] = !f[712] && f[370] && !f[286] && f[492];
	assign leaf[7662] = !f[712] && f[370] && f[286] && !f[316];
	assign leaf[7663] = !f[712] && f[370] && f[286] && f[316];
	assign leaf[7664] = f[712] && !f[231] && !f[295] && !f[689];
	assign leaf[7665] = f[712] && !f[231] && !f[295] && f[689];
	assign leaf[7666] = f[712] && !f[231] && f[295] && !f[180];
	assign leaf[7667] = f[712] && !f[231] && f[295] && f[180];
	assign leaf[7668] = f[712] && f[231] && !f[465] && !f[604];
	assign leaf[7669] = f[712] && f[231] && !f[465] && f[604];
	assign leaf[7670] = f[712] && f[231] && f[465] && !f[578];
	assign leaf[7671] = f[712] && f[231] && f[465] && f[578];
	
	// Tree 544, Classifier 4, Iteration: 54
	assign leaf[7672] = !f[72] && !f[741] && !f[94] && !f[737];
	assign leaf[7673] = !f[72] && !f[741] && !f[94] && f[737];
	assign leaf[7674] = !f[72] && !f[741] && f[94];
	assign leaf[7675] = !f[72] && f[741] && !f[264] && !f[321];
	assign leaf[7676] = !f[72] && f[741] && !f[264] && f[321];
	assign leaf[7677] = !f[72] && f[741] && f[264];
	assign leaf[7678] = f[72];
	
	// Tree 545, Classifier 5, Iteration: 54
	assign leaf[7679] = !f[382] && !f[440] && !f[324] && !f[270];
	assign leaf[7680] = !f[382] && !f[440] && !f[324] && f[270];
	assign leaf[7681] = !f[382] && !f[440] && f[324] && !f[328];
	assign leaf[7682] = !f[382] && !f[440] && f[324] && f[328];
	assign leaf[7683] = !f[382] && f[440] && !f[327] && !f[582];
	assign leaf[7684] = !f[382] && f[440] && !f[327] && f[582];
	assign leaf[7685] = !f[382] && f[440] && f[327] && !f[272];
	assign leaf[7686] = !f[382] && f[440] && f[327] && f[272];
	assign leaf[7687] = f[382] && !f[328] && !f[464] && !f[217];
	assign leaf[7688] = f[382] && !f[328] && !f[464] && f[217];
	assign leaf[7689] = f[382] && !f[328] && f[464] && !f[323];
	assign leaf[7690] = f[382] && !f[328] && f[464] && f[323];
	assign leaf[7691] = f[382] && f[328] && !f[324] && !f[636];
	assign leaf[7692] = f[382] && f[328] && !f[324] && f[636];
	assign leaf[7693] = f[382] && f[328] && f[324] && !f[272];
	assign leaf[7694] = f[382] && f[328] && f[324] && f[272];
	
	// Tree 546, Classifier 6, Iteration: 54
	assign leaf[7695] = !f[295] && !f[214] && !f[635] && !f[627];
	assign leaf[7696] = !f[295] && !f[214] && !f[635] && f[627];
	assign leaf[7697] = !f[295] && !f[214] && f[635] && !f[130];
	assign leaf[7698] = !f[295] && !f[214] && f[635] && f[130];
	assign leaf[7699] = !f[295] && f[214] && !f[663] && !f[657];
	assign leaf[7700] = !f[295] && f[214] && !f[663] && f[657];
	assign leaf[7701] = !f[295] && f[214] && f[663];
	assign leaf[7702] = f[295] && !f[237] && !f[291] && !f[321];
	assign leaf[7703] = f[295] && !f[237] && !f[291] && f[321];
	assign leaf[7704] = f[295] && !f[237] && f[291] && !f[207];
	assign leaf[7705] = f[295] && !f[237] && f[291] && f[207];
	assign leaf[7706] = f[295] && f[237] && !f[374] && !f[323];
	assign leaf[7707] = f[295] && f[237] && !f[374] && f[323];
	assign leaf[7708] = f[295] && f[237] && f[374] && !f[155];
	assign leaf[7709] = f[295] && f[237] && f[374] && f[155];
	
	// Tree 547, Classifier 7, Iteration: 54
	assign leaf[7710] = !f[678] && !f[596] && !f[434] && !f[488];
	assign leaf[7711] = !f[678] && !f[596] && !f[434] && f[488];
	assign leaf[7712] = !f[678] && !f[596] && f[434] && !f[490];
	assign leaf[7713] = !f[678] && !f[596] && f[434] && f[490];
	assign leaf[7714] = !f[678] && f[596] && !f[542] && !f[399];
	assign leaf[7715] = !f[678] && f[596] && !f[542] && f[399];
	assign leaf[7716] = !f[678] && f[596] && f[542] && !f[546];
	assign leaf[7717] = !f[678] && f[596] && f[542] && f[546];
	assign leaf[7718] = f[678] && !f[597] && !f[325];
	assign leaf[7719] = f[678] && !f[597] && f[325];
	assign leaf[7720] = f[678] && f[597] && !f[521] && !f[404];
	assign leaf[7721] = f[678] && f[597] && !f[521] && f[404];
	assign leaf[7722] = f[678] && f[597] && f[521];
	
	// Tree 548, Classifier 8, Iteration: 54
	assign leaf[7723] = !f[176] && !f[687] && !f[630] && !f[575];
	assign leaf[7724] = !f[176] && !f[687] && !f[630] && f[575];
	assign leaf[7725] = !f[176] && !f[687] && f[630] && !f[657];
	assign leaf[7726] = !f[176] && !f[687] && f[630] && f[657];
	assign leaf[7727] = !f[176] && f[687] && !f[631] && !f[689];
	assign leaf[7728] = !f[176] && f[687] && !f[631] && f[689];
	assign leaf[7729] = !f[176] && f[687] && f[631] && !f[545];
	assign leaf[7730] = !f[176] && f[687] && f[631] && f[545];
	assign leaf[7731] = f[176] && !f[657] && !f[636] && !f[628];
	assign leaf[7732] = f[176] && !f[657] && !f[636] && f[628];
	assign leaf[7733] = f[176] && !f[657] && f[636] && !f[631];
	assign leaf[7734] = f[176] && !f[657] && f[636] && f[631];
	assign leaf[7735] = f[176] && f[657] && !f[209] && !f[128];
	assign leaf[7736] = f[176] && f[657] && !f[209] && f[128];
	assign leaf[7737] = f[176] && f[657] && f[209] && !f[492];
	assign leaf[7738] = f[176] && f[657] && f[209] && f[492];
	
	// Tree 549, Classifier 9, Iteration: 54
	assign leaf[7739] = !f[323] && !f[355] && !f[297] && !f[463];
	assign leaf[7740] = !f[323] && !f[355] && !f[297] && f[463];
	assign leaf[7741] = !f[323] && !f[355] && f[297] && !f[241];
	assign leaf[7742] = !f[323] && !f[355] && f[297] && f[241];
	assign leaf[7743] = !f[323] && f[355] && !f[407] && !f[515];
	assign leaf[7744] = !f[323] && f[355] && !f[407] && f[515];
	assign leaf[7745] = !f[323] && f[355] && f[407] && !f[213];
	assign leaf[7746] = !f[323] && f[355] && f[407] && f[213];
	assign leaf[7747] = f[323] && !f[295] && !f[188] && !f[519];
	assign leaf[7748] = f[323] && !f[295] && !f[188] && f[519];
	assign leaf[7749] = f[323] && !f[295] && f[188] && !f[683];
	assign leaf[7750] = f[323] && !f[295] && f[188] && f[683];
	assign leaf[7751] = f[323] && f[295] && !f[575] && !f[179];
	assign leaf[7752] = f[323] && f[295] && !f[575] && f[179];
	assign leaf[7753] = f[323] && f[295] && f[575] && !f[489];
	assign leaf[7754] = f[323] && f[295] && f[575] && f[489];
	
	// Tree 550, Classifier 0, Iteration: 55
	assign leaf[7755] = !f[444] && !f[609] && !f[402] && !f[494];
	assign leaf[7756] = !f[444] && !f[609] && !f[402] && f[494];
	assign leaf[7757] = !f[444] && !f[609] && f[402] && !f[347];
	assign leaf[7758] = !f[444] && !f[609] && f[402] && f[347];
	assign leaf[7759] = !f[444] && f[609] && !f[180] && !f[232];
	assign leaf[7760] = !f[444] && f[609] && !f[180] && f[232];
	assign leaf[7761] = !f[444] && f[609] && f[180] && !f[347];
	assign leaf[7762] = !f[444] && f[609] && f[180] && f[347];
	assign leaf[7763] = f[444] && !f[152] && !f[317];
	assign leaf[7764] = f[444] && !f[152] && f[317] && !f[359];
	assign leaf[7765] = f[444] && !f[152] && f[317] && f[359];
	assign leaf[7766] = f[444] && f[152] && !f[272];
	assign leaf[7767] = f[444] && f[152] && f[272];
	
	// Tree 551, Classifier 1, Iteration: 55
	assign leaf[7768] = !f[683] && !f[411] && !f[556] && !f[606];
	assign leaf[7769] = !f[683] && !f[411] && !f[556] && f[606];
	assign leaf[7770] = !f[683] && !f[411] && f[556];
	assign leaf[7771] = !f[683] && f[411] && !f[156];
	assign leaf[7772] = !f[683] && f[411] && f[156];
	assign leaf[7773] = f[683] && !f[268];
	assign leaf[7774] = f[683] && f[268] && !f[207] && !f[352];
	assign leaf[7775] = f[683] && f[268] && !f[207] && f[352];
	assign leaf[7776] = f[683] && f[268] && f[207];
	
	// Tree 552, Classifier 2, Iteration: 55
	assign leaf[7777] = !f[378] && !f[400] && !f[425] && !f[149];
	assign leaf[7778] = !f[378] && !f[400] && !f[425] && f[149];
	assign leaf[7779] = !f[378] && !f[400] && f[425] && !f[433];
	assign leaf[7780] = !f[378] && !f[400] && f[425] && f[433];
	assign leaf[7781] = !f[378] && f[400] && !f[404] && !f[456];
	assign leaf[7782] = !f[378] && f[400] && !f[404] && f[456];
	assign leaf[7783] = !f[378] && f[400] && f[404] && !f[343];
	assign leaf[7784] = !f[378] && f[400] && f[404] && f[343];
	assign leaf[7785] = f[378] && !f[484] && !f[516] && !f[426];
	assign leaf[7786] = f[378] && !f[484] && !f[516] && f[426];
	assign leaf[7787] = f[378] && !f[484] && f[516] && !f[579];
	assign leaf[7788] = f[378] && !f[484] && f[516] && f[579];
	assign leaf[7789] = f[378] && f[484] && !f[690] && !f[314];
	assign leaf[7790] = f[378] && f[484] && !f[690] && f[314];
	assign leaf[7791] = f[378] && f[484] && f[690];
	
	// Tree 553, Classifier 3, Iteration: 55
	assign leaf[7792] = !f[241] && !f[203] && !f[147] && !f[244];
	assign leaf[7793] = !f[241] && !f[203] && !f[147] && f[244];
	assign leaf[7794] = !f[241] && !f[203] && f[147] && !f[264];
	assign leaf[7795] = !f[241] && !f[203] && f[147] && f[264];
	assign leaf[7796] = !f[241] && f[203] && !f[259] && !f[492];
	assign leaf[7797] = !f[241] && f[203] && !f[259] && f[492];
	assign leaf[7798] = !f[241] && f[203] && f[259] && !f[434];
	assign leaf[7799] = !f[241] && f[203] && f[259] && f[434];
	assign leaf[7800] = f[241] && !f[347] && !f[290] && !f[372];
	assign leaf[7801] = f[241] && !f[347] && !f[290] && f[372];
	assign leaf[7802] = f[241] && !f[347] && f[290] && !f[179];
	assign leaf[7803] = f[241] && !f[347] && f[290] && f[179];
	assign leaf[7804] = f[241] && f[347] && !f[264] && !f[289];
	assign leaf[7805] = f[241] && f[347] && !f[264] && f[289];
	assign leaf[7806] = f[241] && f[347] && f[264] && !f[295];
	assign leaf[7807] = f[241] && f[347] && f[264] && f[295];
	
	// Tree 554, Classifier 4, Iteration: 55
	assign leaf[7808] = !f[318] && !f[320] && !f[316] && !f[230];
	assign leaf[7809] = !f[318] && !f[320] && !f[316] && f[230];
	assign leaf[7810] = !f[318] && !f[320] && f[316] && !f[181];
	assign leaf[7811] = !f[318] && !f[320] && f[316] && f[181];
	assign leaf[7812] = !f[318] && f[320] && !f[262] && !f[347];
	assign leaf[7813] = !f[318] && f[320] && !f[262] && f[347];
	assign leaf[7814] = !f[318] && f[320] && f[262] && !f[633];
	assign leaf[7815] = !f[318] && f[320] && f[262] && f[633];
	assign leaf[7816] = f[318] && !f[321] && !f[209] && !f[265];
	assign leaf[7817] = f[318] && !f[321] && !f[209] && f[265];
	assign leaf[7818] = f[318] && !f[321] && f[209] && !f[212];
	assign leaf[7819] = f[318] && !f[321] && f[209] && f[212];
	assign leaf[7820] = f[318] && f[321] && !f[289] && !f[401];
	assign leaf[7821] = f[318] && f[321] && !f[289] && f[401];
	assign leaf[7822] = f[318] && f[321] && f[289] && !f[291];
	assign leaf[7823] = f[318] && f[321] && f[289] && f[291];
	
	// Tree 555, Classifier 5, Iteration: 55
	assign leaf[7824] = !f[583] && !f[386] && !f[471] && !f[331];
	assign leaf[7825] = !f[583] && !f[386] && !f[471] && f[331];
	assign leaf[7826] = !f[583] && !f[386] && f[471] && !f[354];
	assign leaf[7827] = !f[583] && !f[386] && f[471] && f[354];
	assign leaf[7828] = !f[583] && f[386] && !f[302] && !f[658];
	assign leaf[7829] = !f[583] && f[386] && !f[302] && f[658];
	assign leaf[7830] = !f[583] && f[386] && f[302];
	assign leaf[7831] = f[583] && !f[230] && !f[176] && !f[398];
	assign leaf[7832] = f[583] && !f[230] && !f[176] && f[398];
	assign leaf[7833] = f[583] && !f[230] && f[176] && !f[408];
	assign leaf[7834] = f[583] && !f[230] && f[176] && f[408];
	assign leaf[7835] = f[583] && f[230] && !f[287];
	assign leaf[7836] = f[583] && f[230] && f[287] && !f[238];
	assign leaf[7837] = f[583] && f[230] && f[287] && f[238];
	
	// Tree 556, Classifier 6, Iteration: 55
	assign leaf[7838] = !f[639] && !f[517] && !f[512] && !f[407];
	assign leaf[7839] = !f[639] && !f[517] && !f[512] && f[407];
	assign leaf[7840] = !f[639] && !f[517] && f[512] && !f[373];
	assign leaf[7841] = !f[639] && !f[517] && f[512] && f[373];
	assign leaf[7842] = !f[639] && f[517] && !f[574] && !f[515];
	assign leaf[7843] = !f[639] && f[517] && !f[574] && f[515];
	assign leaf[7844] = !f[639] && f[517] && f[574] && !f[239];
	assign leaf[7845] = !f[639] && f[517] && f[574] && f[239];
	assign leaf[7846] = f[639];
	
	// Tree 557, Classifier 7, Iteration: 55
	assign leaf[7847] = !f[122] && !f[148] && !f[160] && !f[600];
	assign leaf[7848] = !f[122] && !f[148] && !f[160] && f[600];
	assign leaf[7849] = !f[122] && !f[148] && f[160] && !f[651];
	assign leaf[7850] = !f[122] && !f[148] && f[160] && f[651];
	assign leaf[7851] = !f[122] && f[148] && !f[153] && !f[173];
	assign leaf[7852] = !f[122] && f[148] && !f[153] && f[173];
	assign leaf[7853] = !f[122] && f[148] && f[153] && !f[548];
	assign leaf[7854] = !f[122] && f[148] && f[153] && f[548];
	assign leaf[7855] = f[122];
	
	// Tree 558, Classifier 8, Iteration: 55
	assign leaf[7856] = !f[525] && !f[570] && !f[540] && !f[572];
	assign leaf[7857] = !f[525] && !f[570] && !f[540] && f[572];
	assign leaf[7858] = !f[525] && !f[570] && f[540] && !f[604];
	assign leaf[7859] = !f[525] && !f[570] && f[540] && f[604];
	assign leaf[7860] = !f[525] && f[570] && !f[572] && !f[518];
	assign leaf[7861] = !f[525] && f[570] && !f[572] && f[518];
	assign leaf[7862] = !f[525] && f[570] && f[572] && !f[296];
	assign leaf[7863] = !f[525] && f[570] && f[572] && f[296];
	assign leaf[7864] = f[525] && !f[470] && !f[296] && !f[523];
	assign leaf[7865] = f[525] && !f[470] && !f[296] && f[523];
	assign leaf[7866] = f[525] && !f[470] && f[296] && !f[550];
	assign leaf[7867] = f[525] && !f[470] && f[296] && f[550];
	assign leaf[7868] = f[525] && f[470] && !f[456] && !f[438];
	assign leaf[7869] = f[525] && f[470] && !f[456] && f[438];
	assign leaf[7870] = f[525] && f[470] && f[456] && !f[125];
	assign leaf[7871] = f[525] && f[470] && f[456] && f[125];
	
	// Tree 559, Classifier 9, Iteration: 55
	assign leaf[7872] = !f[742] && !f[686] && !f[740] && !f[602];
	assign leaf[7873] = !f[742] && !f[686] && !f[740] && f[602];
	assign leaf[7874] = !f[742] && !f[686] && f[740] && !f[710];
	assign leaf[7875] = !f[742] && !f[686] && f[740] && f[710];
	assign leaf[7876] = !f[742] && f[686] && !f[545] && !f[408];
	assign leaf[7877] = !f[742] && f[686] && !f[545] && f[408];
	assign leaf[7878] = !f[742] && f[686] && f[545] && !f[184];
	assign leaf[7879] = !f[742] && f[686] && f[545] && f[184];
	assign leaf[7880] = f[742] && !f[242] && !f[405] && !f[322];
	assign leaf[7881] = f[742] && !f[242] && !f[405] && f[322];
	assign leaf[7882] = f[742] && !f[242] && f[405] && !f[326];
	assign leaf[7883] = f[742] && !f[242] && f[405] && f[326];
	assign leaf[7884] = f[742] && f[242] && !f[684] && !f[488];
	assign leaf[7885] = f[742] && f[242] && !f[684] && f[488];
	assign leaf[7886] = f[742] && f[242] && f[684];
	
	// Tree 560, Classifier 0, Iteration: 56
	assign leaf[7887] = !f[416] && !f[214] && !f[241] && !f[438];
	assign leaf[7888] = !f[416] && !f[214] && !f[241] && f[438];
	assign leaf[7889] = !f[416] && !f[214] && f[241] && !f[542];
	assign leaf[7890] = !f[416] && !f[214] && f[241] && f[542];
	assign leaf[7891] = !f[416] && f[214] && !f[516] && !f[380];
	assign leaf[7892] = !f[416] && f[214] && !f[516] && f[380];
	assign leaf[7893] = !f[416] && f[214] && f[516] && !f[186];
	assign leaf[7894] = !f[416] && f[214] && f[516] && f[186];
	assign leaf[7895] = f[416] && !f[398];
	assign leaf[7896] = f[416] && f[398] && !f[289];
	assign leaf[7897] = f[416] && f[398] && f[289] && !f[430];
	assign leaf[7898] = f[416] && f[398] && f[289] && f[430];
	
	// Tree 561, Classifier 1, Iteration: 56
	assign leaf[7899] = !f[583] && !f[152] && !f[98] && !f[236];
	assign leaf[7900] = !f[583] && !f[152] && !f[98] && f[236];
	assign leaf[7901] = !f[583] && !f[152] && f[98] && !f[236];
	assign leaf[7902] = !f[583] && !f[152] && f[98] && f[236];
	assign leaf[7903] = !f[583] && f[152] && !f[269] && !f[265];
	assign leaf[7904] = !f[583] && f[152] && !f[269] && f[265];
	assign leaf[7905] = !f[583] && f[152] && f[269] && !f[604];
	assign leaf[7906] = !f[583] && f[152] && f[269] && f[604];
	assign leaf[7907] = f[583];
	
	// Tree 562, Classifier 2, Iteration: 56
	assign leaf[7908] = !f[418] && !f[411] && !f[329] && !f[378];
	assign leaf[7909] = !f[418] && !f[411] && !f[329] && f[378];
	assign leaf[7910] = !f[418] && !f[411] && f[329] && !f[324];
	assign leaf[7911] = !f[418] && !f[411] && f[329] && f[324];
	assign leaf[7912] = !f[418] && f[411] && !f[353] && !f[540];
	assign leaf[7913] = !f[418] && f[411] && !f[353] && f[540];
	assign leaf[7914] = !f[418] && f[411] && f[353] && !f[519];
	assign leaf[7915] = !f[418] && f[411] && f[353] && f[519];
	assign leaf[7916] = f[418];
	
	// Tree 563, Classifier 3, Iteration: 56
	assign leaf[7917] = !f[369] && !f[402] && !f[544] && !f[211];
	assign leaf[7918] = !f[369] && !f[402] && !f[544] && f[211];
	assign leaf[7919] = !f[369] && !f[402] && f[544] && !f[547];
	assign leaf[7920] = !f[369] && !f[402] && f[544] && f[547];
	assign leaf[7921] = !f[369] && f[402] && !f[526] && !f[318];
	assign leaf[7922] = !f[369] && f[402] && !f[526] && f[318];
	assign leaf[7923] = !f[369] && f[402] && f[526] && !f[126];
	assign leaf[7924] = !f[369] && f[402] && f[526] && f[126];
	assign leaf[7925] = f[369] && !f[544] && !f[217] && !f[293];
	assign leaf[7926] = f[369] && !f[544] && !f[217] && f[293];
	assign leaf[7927] = f[369] && !f[544] && f[217];
	assign leaf[7928] = f[369] && f[544] && !f[234];
	assign leaf[7929] = f[369] && f[544] && f[234];
	
	// Tree 564, Classifier 4, Iteration: 56
	assign leaf[7930] = !f[430] && !f[569] && !f[549] && !f[413];
	assign leaf[7931] = !f[430] && !f[569] && !f[549] && f[413];
	assign leaf[7932] = !f[430] && !f[569] && f[549] && !f[691];
	assign leaf[7933] = !f[430] && !f[569] && f[549] && f[691];
	assign leaf[7934] = !f[430] && f[569] && !f[497] && !f[680];
	assign leaf[7935] = !f[430] && f[569] && !f[497] && f[680];
	assign leaf[7936] = !f[430] && f[569] && f[497];
	assign leaf[7937] = f[430] && !f[206] && !f[662] && !f[152];
	assign leaf[7938] = f[430] && !f[206] && !f[662] && f[152];
	assign leaf[7939] = f[430] && !f[206] && f[662] && !f[659];
	assign leaf[7940] = f[430] && !f[206] && f[662] && f[659];
	assign leaf[7941] = f[430] && f[206] && !f[237] && !f[155];
	assign leaf[7942] = f[430] && f[206] && !f[237] && f[155];
	assign leaf[7943] = f[430] && f[206] && f[237] && !f[272];
	assign leaf[7944] = f[430] && f[206] && f[237] && f[272];
	
	// Tree 565, Classifier 5, Iteration: 56
	assign leaf[7945] = !f[598] && !f[214] && !f[270] && !f[266];
	assign leaf[7946] = !f[598] && !f[214] && !f[270] && f[266];
	assign leaf[7947] = !f[598] && !f[214] && f[270] && !f[294];
	assign leaf[7948] = !f[598] && !f[214] && f[270] && f[294];
	assign leaf[7949] = !f[598] && f[214] && !f[297] && !f[327];
	assign leaf[7950] = !f[598] && f[214] && !f[297] && f[327];
	assign leaf[7951] = !f[598] && f[214] && f[297] && !f[709];
	assign leaf[7952] = !f[598] && f[214] && f[297] && f[709];
	assign leaf[7953] = f[598] && !f[486] && !f[428] && !f[398];
	assign leaf[7954] = f[598] && !f[486] && !f[428] && f[398];
	assign leaf[7955] = f[598] && !f[486] && f[428] && !f[483];
	assign leaf[7956] = f[598] && !f[486] && f[428] && f[483];
	assign leaf[7957] = f[598] && f[486] && !f[541] && !f[429];
	assign leaf[7958] = f[598] && f[486] && !f[541] && f[429];
	assign leaf[7959] = f[598] && f[486] && f[541] && !f[370];
	assign leaf[7960] = f[598] && f[486] && f[541] && f[370];
	
	// Tree 566, Classifier 6, Iteration: 56
	assign leaf[7961] = !f[684] && !f[302] && !f[455] && !f[288];
	assign leaf[7962] = !f[684] && !f[302] && !f[455] && f[288];
	assign leaf[7963] = !f[684] && !f[302] && f[455] && !f[511];
	assign leaf[7964] = !f[684] && !f[302] && f[455] && f[511];
	assign leaf[7965] = !f[684] && f[302] && !f[402] && !f[298];
	assign leaf[7966] = !f[684] && f[302] && !f[402] && f[298];
	assign leaf[7967] = !f[684] && f[302] && f[402] && !f[127];
	assign leaf[7968] = !f[684] && f[302] && f[402] && f[127];
	assign leaf[7969] = f[684] && !f[513];
	assign leaf[7970] = f[684] && f[513];
	
	// Tree 567, Classifier 7, Iteration: 56
	assign leaf[7971] = !f[583] && !f[122] && !f[183] && !f[488];
	assign leaf[7972] = !f[583] && !f[122] && !f[183] && f[488];
	assign leaf[7973] = !f[583] && !f[122] && f[183] && !f[320];
	assign leaf[7974] = !f[583] && !f[122] && f[183] && f[320];
	assign leaf[7975] = !f[583] && f[122];
	assign leaf[7976] = f[583];
	
	// Tree 568, Classifier 8, Iteration: 56
	assign leaf[7977] = !f[341] && !f[277] && !f[679] && !f[302];
	assign leaf[7978] = !f[341] && !f[277] && !f[679] && f[302];
	assign leaf[7979] = !f[341] && !f[277] && f[679] && !f[540];
	assign leaf[7980] = !f[341] && !f[277] && f[679] && f[540];
	assign leaf[7981] = !f[341] && f[277] && !f[401];
	assign leaf[7982] = !f[341] && f[277] && f[401] && !f[383];
	assign leaf[7983] = !f[341] && f[277] && f[401] && f[383];
	assign leaf[7984] = f[341] && !f[315] && !f[625] && !f[177];
	assign leaf[7985] = f[341] && !f[315] && !f[625] && f[177];
	assign leaf[7986] = f[341] && !f[315] && f[625];
	assign leaf[7987] = f[341] && f[315] && !f[264] && !f[572];
	assign leaf[7988] = f[341] && f[315] && !f[264] && f[572];
	assign leaf[7989] = f[341] && f[315] && f[264] && !f[383];
	assign leaf[7990] = f[341] && f[315] && f[264] && f[383];
	
	// Tree 569, Classifier 9, Iteration: 56
	assign leaf[7991] = !f[131] && !f[369] && !f[441] && !f[497];
	assign leaf[7992] = !f[131] && !f[369] && !f[441] && f[497];
	assign leaf[7993] = !f[131] && !f[369] && f[441] && !f[544];
	assign leaf[7994] = !f[131] && !f[369] && f[441] && f[544];
	assign leaf[7995] = !f[131] && f[369] && !f[346] && !f[359];
	assign leaf[7996] = !f[131] && f[369] && !f[346] && f[359];
	assign leaf[7997] = !f[131] && f[369] && f[346] && !f[386];
	assign leaf[7998] = !f[131] && f[369] && f[346] && f[386];
	assign leaf[7999] = f[131] && !f[509];
	assign leaf[8000] = f[131] && f[509];
	
	// Tree 570, Classifier 0, Iteration: 57
	assign leaf[8001] = !f[434] && !f[664] && !f[433] && !f[547];
	assign leaf[8002] = !f[434] && !f[664] && !f[433] && f[547];
	assign leaf[8003] = !f[434] && !f[664] && f[433] && !f[348];
	assign leaf[8004] = !f[434] && !f[664] && f[433] && f[348];
	assign leaf[8005] = !f[434] && f[664] && !f[151];
	assign leaf[8006] = !f[434] && f[664] && f[151];
	assign leaf[8007] = f[434] && !f[456] && !f[386];
	assign leaf[8008] = f[434] && !f[456] && f[386];
	assign leaf[8009] = f[434] && f[456] && !f[461] && !f[267];
	assign leaf[8010] = f[434] && f[456] && !f[461] && f[267];
	assign leaf[8011] = f[434] && f[456] && f[461] && !f[357];
	assign leaf[8012] = f[434] && f[456] && f[461] && f[357];
	
	// Tree 571, Classifier 1, Iteration: 57
	assign leaf[8013] = !f[604] && !f[180] && !f[320] && !f[492];
	assign leaf[8014] = !f[604] && !f[180] && !f[320] && f[492];
	assign leaf[8015] = !f[604] && !f[180] && f[320] && !f[631];
	assign leaf[8016] = !f[604] && !f[180] && f[320] && f[631];
	assign leaf[8017] = !f[604] && f[180] && !f[269] && !f[236];
	assign leaf[8018] = !f[604] && f[180] && !f[269] && f[236];
	assign leaf[8019] = !f[604] && f[180] && f[269] && !f[207];
	assign leaf[8020] = !f[604] && f[180] && f[269] && f[207];
	assign leaf[8021] = f[604] && !f[547] && !f[266] && !f[569];
	assign leaf[8022] = f[604] && !f[547] && !f[266] && f[569];
	assign leaf[8023] = f[604] && !f[547] && f[266] && !f[493];
	assign leaf[8024] = f[604] && !f[547] && f[266] && f[493];
	assign leaf[8025] = f[604] && f[547] && !f[488] && !f[350];
	assign leaf[8026] = f[604] && f[547] && !f[488] && f[350];
	assign leaf[8027] = f[604] && f[547] && f[488] && !f[574];
	assign leaf[8028] = f[604] && f[547] && f[488] && f[574];
	
	// Tree 572, Classifier 2, Iteration: 57
	assign leaf[8029] = !f[513] && !f[404] && !f[568] && !f[458];
	assign leaf[8030] = !f[513] && !f[404] && !f[568] && f[458];
	assign leaf[8031] = !f[513] && !f[404] && f[568] && !f[320];
	assign leaf[8032] = !f[513] && !f[404] && f[568] && f[320];
	assign leaf[8033] = !f[513] && f[404] && !f[455] && !f[97];
	assign leaf[8034] = !f[513] && f[404] && !f[455] && f[97];
	assign leaf[8035] = !f[513] && f[404] && f[455] && !f[401];
	assign leaf[8036] = !f[513] && f[404] && f[455] && f[401];
	assign leaf[8037] = f[513] && !f[459] && !f[351] && !f[552];
	assign leaf[8038] = f[513] && !f[459] && !f[351] && f[552];
	assign leaf[8039] = f[513] && !f[459] && f[351] && !f[430];
	assign leaf[8040] = f[513] && !f[459] && f[351] && f[430];
	assign leaf[8041] = f[513] && f[459] && !f[294] && !f[186];
	assign leaf[8042] = f[513] && f[459] && !f[294] && f[186];
	assign leaf[8043] = f[513] && f[459] && f[294] && !f[96];
	assign leaf[8044] = f[513] && f[459] && f[294] && f[96];
	
	// Tree 573, Classifier 3, Iteration: 57
	assign leaf[8045] = !f[708] && !f[357] && !f[190] && !f[649];
	assign leaf[8046] = !f[708] && !f[357] && !f[190] && f[649];
	assign leaf[8047] = !f[708] && !f[357] && f[190] && !f[355];
	assign leaf[8048] = !f[708] && !f[357] && f[190] && f[355];
	assign leaf[8049] = !f[708] && f[357] && !f[266] && !f[160];
	assign leaf[8050] = !f[708] && f[357] && !f[266] && f[160];
	assign leaf[8051] = !f[708] && f[357] && f[266] && !f[187];
	assign leaf[8052] = !f[708] && f[357] && f[266] && f[187];
	assign leaf[8053] = f[708] && !f[599] && !f[518] && !f[244];
	assign leaf[8054] = f[708] && !f[599] && !f[518] && f[244];
	assign leaf[8055] = f[708] && !f[599] && f[518];
	assign leaf[8056] = f[708] && f[599] && !f[602];
	assign leaf[8057] = f[708] && f[599] && f[602];
	
	// Tree 574, Classifier 4, Iteration: 57
	assign leaf[8058] = !f[430] && !f[300] && !f[181] && !f[265];
	assign leaf[8059] = !f[430] && !f[300] && !f[181] && f[265];
	assign leaf[8060] = !f[430] && !f[300] && f[181] && !f[234];
	assign leaf[8061] = !f[430] && !f[300] && f[181] && f[234];
	assign leaf[8062] = !f[430] && f[300] && !f[182] && !f[206];
	assign leaf[8063] = !f[430] && f[300] && !f[182] && f[206];
	assign leaf[8064] = !f[430] && f[300] && f[182] && !f[185];
	assign leaf[8065] = !f[430] && f[300] && f[182] && f[185];
	assign leaf[8066] = f[430] && !f[427] && !f[581] && !f[626];
	assign leaf[8067] = f[430] && !f[427] && !f[581] && f[626];
	assign leaf[8068] = f[430] && !f[427] && f[581] && !f[353];
	assign leaf[8069] = f[430] && !f[427] && f[581] && f[353];
	assign leaf[8070] = f[430] && f[427] && !f[513] && !f[435];
	assign leaf[8071] = f[430] && f[427] && !f[513] && f[435];
	assign leaf[8072] = f[430] && f[427] && f[513] && !f[497];
	assign leaf[8073] = f[430] && f[427] && f[513] && f[497];
	
	// Tree 575, Classifier 5, Iteration: 57
	assign leaf[8074] = !f[129] && !f[215] && !f[273] && !f[239];
	assign leaf[8075] = !f[129] && !f[215] && !f[273] && f[239];
	assign leaf[8076] = !f[129] && !f[215] && f[273] && !f[270];
	assign leaf[8077] = !f[129] && !f[215] && f[273] && f[270];
	assign leaf[8078] = !f[129] && f[215] && !f[297] && !f[328];
	assign leaf[8079] = !f[129] && f[215] && !f[297] && f[328];
	assign leaf[8080] = !f[129] && f[215] && f[297] && !f[293];
	assign leaf[8081] = !f[129] && f[215] && f[297] && f[293];
	assign leaf[8082] = f[129] && !f[242] && !f[218] && !f[601];
	assign leaf[8083] = f[129] && !f[242] && !f[218] && f[601];
	assign leaf[8084] = f[129] && !f[242] && f[218];
	assign leaf[8085] = f[129] && f[242] && !f[239];
	assign leaf[8086] = f[129] && f[242] && f[239] && !f[125];
	assign leaf[8087] = f[129] && f[242] && f[239] && f[125];
	
	// Tree 576, Classifier 6, Iteration: 57
	assign leaf[8088] = !f[495] && !f[494] && !f[497] && !f[131];
	assign leaf[8089] = !f[495] && !f[494] && !f[497] && f[131];
	assign leaf[8090] = !f[495] && !f[494] && f[497] && !f[348];
	assign leaf[8091] = !f[495] && !f[494] && f[497] && f[348];
	assign leaf[8092] = !f[495] && f[494] && !f[234] && !f[544];
	assign leaf[8093] = !f[495] && f[494] && !f[234] && f[544];
	assign leaf[8094] = !f[495] && f[494] && f[234] && !f[439];
	assign leaf[8095] = !f[495] && f[494] && f[234] && f[439];
	assign leaf[8096] = f[495] && !f[431] && !f[464] && !f[434];
	assign leaf[8097] = f[495] && !f[431] && !f[464] && f[434];
	assign leaf[8098] = f[495] && !f[431] && f[464] && !f[487];
	assign leaf[8099] = f[495] && !f[431] && f[464] && f[487];
	assign leaf[8100] = f[495] && f[431] && !f[230] && !f[302];
	assign leaf[8101] = f[495] && f[431] && !f[230] && f[302];
	assign leaf[8102] = f[495] && f[431] && f[230];
	
	// Tree 577, Classifier 7, Iteration: 57
	assign leaf[8103] = !f[359] && !f[202] && !f[548] && !f[603];
	assign leaf[8104] = !f[359] && !f[202] && !f[548] && f[603];
	assign leaf[8105] = !f[359] && !f[202] && f[548] && !f[433];
	assign leaf[8106] = !f[359] && !f[202] && f[548] && f[433];
	assign leaf[8107] = !f[359] && f[202] && !f[492] && !f[205];
	assign leaf[8108] = !f[359] && f[202] && !f[492] && f[205];
	assign leaf[8109] = !f[359] && f[202] && f[492] && !f[540];
	assign leaf[8110] = !f[359] && f[202] && f[492] && f[540];
	assign leaf[8111] = f[359] && !f[240] && !f[542] && !f[319];
	assign leaf[8112] = f[359] && !f[240] && !f[542] && f[319];
	assign leaf[8113] = f[359] && !f[240] && f[542];
	assign leaf[8114] = f[359] && f[240] && !f[466] && !f[545];
	assign leaf[8115] = f[359] && f[240] && !f[466] && f[545];
	assign leaf[8116] = f[359] && f[240] && f[466] && !f[710];
	assign leaf[8117] = f[359] && f[240] && f[466] && f[710];
	
	// Tree 578, Classifier 8, Iteration: 57
	assign leaf[8118] = !f[165] && !f[381] && !f[464] && !f[491];
	assign leaf[8119] = !f[165] && !f[381] && !f[464] && f[491];
	assign leaf[8120] = !f[165] && !f[381] && f[464] && !f[376];
	assign leaf[8121] = !f[165] && !f[381] && f[464] && f[376];
	assign leaf[8122] = !f[165] && f[381] && !f[297] && !f[295];
	assign leaf[8123] = !f[165] && f[381] && !f[297] && f[295];
	assign leaf[8124] = !f[165] && f[381] && f[297] && !f[180];
	assign leaf[8125] = !f[165] && f[381] && f[297] && f[180];
	assign leaf[8126] = f[165];
	
	// Tree 579, Classifier 9, Iteration: 57
	assign leaf[8127] = !f[734] && !f[380] && !f[440] && !f[325];
	assign leaf[8128] = !f[734] && !f[380] && !f[440] && f[325];
	assign leaf[8129] = !f[734] && !f[380] && f[440] && !f[543];
	assign leaf[8130] = !f[734] && !f[380] && f[440] && f[543];
	assign leaf[8131] = !f[734] && f[380] && !f[467] && !f[523];
	assign leaf[8132] = !f[734] && f[380] && !f[467] && f[523];
	assign leaf[8133] = !f[734] && f[380] && f[467] && !f[343];
	assign leaf[8134] = !f[734] && f[380] && f[467] && f[343];
	assign leaf[8135] = f[734] && !f[597];
	assign leaf[8136] = f[734] && f[597];
	
	// Tree 580, Classifier 0, Iteration: 58
	assign leaf[8137] = !f[688] && !f[663] && !f[712] && !f[397];
	assign leaf[8138] = !f[688] && !f[663] && !f[712] && f[397];
	assign leaf[8139] = !f[688] && !f[663] && f[712] && !f[573];
	assign leaf[8140] = !f[688] && !f[663] && f[712] && f[573];
	assign leaf[8141] = !f[688] && f[663] && !f[659];
	assign leaf[8142] = !f[688] && f[663] && f[659];
	assign leaf[8143] = f[688] && !f[548] && !f[287] && !f[356];
	assign leaf[8144] = f[688] && !f[548] && !f[287] && f[356];
	assign leaf[8145] = f[688] && !f[548] && f[287];
	assign leaf[8146] = f[688] && f[548];
	
	// Tree 581, Classifier 1, Iteration: 58
	assign leaf[8147] = !f[716] && !f[408] && !f[464] && !f[548];
	assign leaf[8148] = !f[716] && !f[408] && !f[464] && f[548];
	assign leaf[8149] = !f[716] && !f[408] && f[464] && !f[268];
	assign leaf[8150] = !f[716] && !f[408] && f[464] && f[268];
	assign leaf[8151] = !f[716] && f[408] && !f[324] && !f[157];
	assign leaf[8152] = !f[716] && f[408] && !f[324] && f[157];
	assign leaf[8153] = !f[716] && f[408] && f[324] && !f[630];
	assign leaf[8154] = !f[716] && f[408] && f[324] && f[630];
	assign leaf[8155] = f[716];
	
	// Tree 582, Classifier 2, Iteration: 58
	assign leaf[8156] = !f[104] && !f[545] && !f[660] && !f[469];
	assign leaf[8157] = !f[104] && !f[545] && !f[660] && f[469];
	assign leaf[8158] = !f[104] && !f[545] && f[660] && !f[464];
	assign leaf[8159] = !f[104] && !f[545] && f[660] && f[464];
	assign leaf[8160] = !f[104] && f[545] && !f[427] && !f[343];
	assign leaf[8161] = !f[104] && f[545] && !f[427] && f[343];
	assign leaf[8162] = !f[104] && f[545] && f[427] && !f[289];
	assign leaf[8163] = !f[104] && f[545] && f[427] && f[289];
	assign leaf[8164] = f[104] && !f[432] && !f[324];
	assign leaf[8165] = f[104] && !f[432] && f[324];
	assign leaf[8166] = f[104] && f[432] && !f[593];
	assign leaf[8167] = f[104] && f[432] && f[593];
	
	// Tree 583, Classifier 3, Iteration: 58
	assign leaf[8168] = !f[384] && !f[495] && !f[293] && !f[298];
	assign leaf[8169] = !f[384] && !f[495] && !f[293] && f[298];
	assign leaf[8170] = !f[384] && !f[495] && f[293] && !f[319];
	assign leaf[8171] = !f[384] && !f[495] && f[293] && f[319];
	assign leaf[8172] = !f[384] && f[495] && !f[442] && !f[435];
	assign leaf[8173] = !f[384] && f[495] && !f[442] && f[435];
	assign leaf[8174] = !f[384] && f[495] && f[442];
	assign leaf[8175] = f[384] && !f[438] && !f[353] && !f[537];
	assign leaf[8176] = f[384] && !f[438] && !f[353] && f[537];
	assign leaf[8177] = f[384] && !f[438] && f[353] && !f[211];
	assign leaf[8178] = f[384] && !f[438] && f[353] && f[211];
	assign leaf[8179] = f[384] && f[438] && !f[517] && !f[327];
	assign leaf[8180] = f[384] && f[438] && !f[517] && f[327];
	assign leaf[8181] = f[384] && f[438] && f[517] && !f[126];
	assign leaf[8182] = f[384] && f[438] && f[517] && f[126];
	
	// Tree 584, Classifier 4, Iteration: 58
	assign leaf[8183] = !f[637] && !f[286] && !f[318] && !f[320];
	assign leaf[8184] = !f[637] && !f[286] && !f[318] && f[320];
	assign leaf[8185] = !f[637] && !f[286] && f[318] && !f[321];
	assign leaf[8186] = !f[637] && !f[286] && f[318] && f[321];
	assign leaf[8187] = !f[637] && f[286] && !f[201] && !f[685];
	assign leaf[8188] = !f[637] && f[286] && !f[201] && f[685];
	assign leaf[8189] = !f[637] && f[286] && f[201];
	assign leaf[8190] = f[637] && !f[234] && !f[151] && !f[523];
	assign leaf[8191] = f[637] && !f[234] && !f[151] && f[523];
	assign leaf[8192] = f[637] && !f[234] && f[151];
	assign leaf[8193] = f[637] && f[234] && !f[482] && !f[462];
	assign leaf[8194] = f[637] && f[234] && !f[482] && f[462];
	assign leaf[8195] = f[637] && f[234] && f[482];
	
	// Tree 585, Classifier 5, Iteration: 58
	assign leaf[8196] = !f[380] && !f[292] && !f[413] && !f[345];
	assign leaf[8197] = !f[380] && !f[292] && !f[413] && f[345];
	assign leaf[8198] = !f[380] && !f[292] && f[413] && !f[661];
	assign leaf[8199] = !f[380] && !f[292] && f[413] && f[661];
	assign leaf[8200] = !f[380] && f[292] && !f[347] && !f[315];
	assign leaf[8201] = !f[380] && f[292] && !f[347] && f[315];
	assign leaf[8202] = !f[380] && f[292] && f[347] && !f[298];
	assign leaf[8203] = !f[380] && f[292] && f[347] && f[298];
	assign leaf[8204] = f[380] && !f[131] && !f[349] && !f[659];
	assign leaf[8205] = f[380] && !f[131] && !f[349] && f[659];
	assign leaf[8206] = f[380] && !f[131] && f[349] && !f[245];
	assign leaf[8207] = f[380] && !f[131] && f[349] && f[245];
	assign leaf[8208] = f[380] && f[131] && !f[630] && !f[550];
	assign leaf[8209] = f[380] && f[131] && !f[630] && f[550];
	assign leaf[8210] = f[380] && f[131] && f[630] && !f[651];
	assign leaf[8211] = f[380] && f[131] && f[630] && f[651];
	
	// Tree 586, Classifier 6, Iteration: 58
	assign leaf[8212] = !f[101] && !f[72] && !f[684] && !f[602];
	assign leaf[8213] = !f[101] && !f[72] && !f[684] && f[602];
	assign leaf[8214] = !f[101] && !f[72] && f[684] && !f[570];
	assign leaf[8215] = !f[101] && !f[72] && f[684] && f[570];
	assign leaf[8216] = !f[101] && f[72];
	assign leaf[8217] = f[101] && !f[293] && !f[521] && !f[209];
	assign leaf[8218] = f[101] && !f[293] && !f[521] && f[209];
	assign leaf[8219] = f[101] && !f[293] && f[521] && !f[463];
	assign leaf[8220] = f[101] && !f[293] && f[521] && f[463];
	assign leaf[8221] = f[101] && f[293] && !f[126] && !f[544];
	assign leaf[8222] = f[101] && f[293] && !f[126] && f[544];
	assign leaf[8223] = f[101] && f[293] && f[126] && !f[626];
	assign leaf[8224] = f[101] && f[293] && f[126] && f[626];
	
	// Tree 587, Classifier 7, Iteration: 58
	assign leaf[8225] = !f[191] && !f[126] && !f[608] && !f[295];
	assign leaf[8226] = !f[191] && !f[126] && !f[608] && f[295];
	assign leaf[8227] = !f[191] && !f[126] && f[608] && !f[270];
	assign leaf[8228] = !f[191] && !f[126] && f[608] && f[270];
	assign leaf[8229] = !f[191] && f[126] && !f[629];
	assign leaf[8230] = !f[191] && f[126] && f[629];
	assign leaf[8231] = f[191] && !f[679];
	assign leaf[8232] = f[191] && f[679];
	
	// Tree 588, Classifier 8, Iteration: 58
	assign leaf[8233] = !f[439] && !f[525] && !f[542] && !f[660];
	assign leaf[8234] = !f[439] && !f[525] && !f[542] && f[660];
	assign leaf[8235] = !f[439] && !f[525] && f[542] && !f[538];
	assign leaf[8236] = !f[439] && !f[525] && f[542] && f[538];
	assign leaf[8237] = !f[439] && f[525] && !f[456] && !f[467];
	assign leaf[8238] = !f[439] && f[525] && !f[456] && f[467];
	assign leaf[8239] = !f[439] && f[525] && f[456] && !f[246];
	assign leaf[8240] = !f[439] && f[525] && f[456] && f[246];
	assign leaf[8241] = f[439] && !f[154] && !f[354] && !f[572];
	assign leaf[8242] = f[439] && !f[154] && !f[354] && f[572];
	assign leaf[8243] = f[439] && !f[154] && f[354] && !f[625];
	assign leaf[8244] = f[439] && !f[154] && f[354] && f[625];
	assign leaf[8245] = f[439] && f[154] && !f[318] && !f[265];
	assign leaf[8246] = f[439] && f[154] && !f[318] && f[265];
	assign leaf[8247] = f[439] && f[154] && f[318] && !f[379];
	assign leaf[8248] = f[439] && f[154] && f[318] && f[379];
	
	// Tree 589, Classifier 9, Iteration: 58
	assign leaf[8249] = !f[149] && !f[388] && !f[508] && !f[256];
	assign leaf[8250] = !f[149] && !f[388] && !f[508] && f[256];
	assign leaf[8251] = !f[149] && !f[388] && f[508] && !f[662];
	assign leaf[8252] = !f[149] && !f[388] && f[508] && f[662];
	assign leaf[8253] = !f[149] && f[388];
	assign leaf[8254] = f[149] && !f[286];
	assign leaf[8255] = f[149] && f[286] && !f[354];
	assign leaf[8256] = f[149] && f[286] && f[354];
	
	// Tree 590, Classifier 0, Iteration: 59
	assign leaf[8257] = !f[380] && !f[512] && !f[271] && !f[403];
	assign leaf[8258] = !f[380] && !f[512] && !f[271] && f[403];
	assign leaf[8259] = !f[380] && !f[512] && f[271] && !f[462];
	assign leaf[8260] = !f[380] && !f[512] && f[271] && f[462];
	assign leaf[8261] = !f[380] && f[512] && !f[429] && !f[359];
	assign leaf[8262] = !f[380] && f[512] && !f[429] && f[359];
	assign leaf[8263] = !f[380] && f[512] && f[429] && !f[353];
	assign leaf[8264] = !f[380] && f[512] && f[429] && f[353];
	assign leaf[8265] = f[380] && !f[268] && !f[314] && !f[126];
	assign leaf[8266] = f[380] && !f[268] && !f[314] && f[126];
	assign leaf[8267] = f[380] && !f[268] && f[314];
	assign leaf[8268] = f[380] && f[268] && !f[325] && !f[329];
	assign leaf[8269] = f[380] && f[268] && !f[325] && f[329];
	assign leaf[8270] = f[380] && f[268] && f[325] && !f[596];
	assign leaf[8271] = f[380] && f[268] && f[325] && f[596];
	
	// Tree 591, Classifier 1, Iteration: 59
	assign leaf[8272] = !f[609] && !f[204] && !f[157] && !f[241];
	assign leaf[8273] = !f[609] && !f[204] && !f[157] && f[241];
	assign leaf[8274] = !f[609] && !f[204] && f[157] && !f[268];
	assign leaf[8275] = !f[609] && !f[204] && f[157] && f[268];
	assign leaf[8276] = !f[609] && f[204] && !f[625] && !f[266];
	assign leaf[8277] = !f[609] && f[204] && !f[625] && f[266];
	assign leaf[8278] = !f[609] && f[204] && f[625];
	assign leaf[8279] = f[609] && !f[157] && !f[548];
	assign leaf[8280] = f[609] && !f[157] && f[548] && !f[516];
	assign leaf[8281] = f[609] && !f[157] && f[548] && f[516];
	assign leaf[8282] = f[609] && f[157];
	
	// Tree 592, Classifier 2, Iteration: 59
	assign leaf[8283] = !f[677] && !f[622] && !f[219] && !f[103];
	assign leaf[8284] = !f[677] && !f[622] && !f[219] && f[103];
	assign leaf[8285] = !f[677] && !f[622] && f[219] && !f[374];
	assign leaf[8286] = !f[677] && !f[622] && f[219] && f[374];
	assign leaf[8287] = !f[677] && f[622] && !f[236] && !f[495];
	assign leaf[8288] = !f[677] && f[622] && !f[236] && f[495];
	assign leaf[8289] = !f[677] && f[622] && f[236] && !f[661];
	assign leaf[8290] = !f[677] && f[622] && f[236] && f[661];
	assign leaf[8291] = f[677] && !f[188];
	assign leaf[8292] = f[677] && f[188];
	
	// Tree 593, Classifier 3, Iteration: 59
	assign leaf[8293] = !f[492] && !f[547] && !f[517] && !f[407];
	assign leaf[8294] = !f[492] && !f[547] && !f[517] && f[407];
	assign leaf[8295] = !f[492] && !f[547] && f[517] && !f[572];
	assign leaf[8296] = !f[492] && !f[547] && f[517] && f[572];
	assign leaf[8297] = !f[492] && f[547] && !f[409] && !f[581];
	assign leaf[8298] = !f[492] && f[547] && !f[409] && f[581];
	assign leaf[8299] = !f[492] && f[547] && f[409] && !f[516];
	assign leaf[8300] = !f[492] && f[547] && f[409] && f[516];
	assign leaf[8301] = f[492] && !f[438] && !f[493] && !f[293];
	assign leaf[8302] = f[492] && !f[438] && !f[493] && f[293];
	assign leaf[8303] = f[492] && !f[438] && f[493] && !f[355];
	assign leaf[8304] = f[492] && !f[438] && f[493] && f[355];
	assign leaf[8305] = f[492] && f[438] && !f[295] && !f[564];
	assign leaf[8306] = f[492] && f[438] && !f[295] && f[564];
	assign leaf[8307] = f[492] && f[438] && f[295] && !f[155];
	assign leaf[8308] = f[492] && f[438] && f[295] && f[155];
	
	// Tree 594, Classifier 4, Iteration: 59
	assign leaf[8309] = !f[743] && !f[398] && !f[347] && !f[181];
	assign leaf[8310] = !f[743] && !f[398] && !f[347] && f[181];
	assign leaf[8311] = !f[743] && !f[398] && f[347] && !f[313];
	assign leaf[8312] = !f[743] && !f[398] && f[347] && f[313];
	assign leaf[8313] = !f[743] && f[398] && !f[344] && !f[343];
	assign leaf[8314] = !f[743] && f[398] && !f[344] && f[343];
	assign leaf[8315] = !f[743] && f[398] && f[344] && !f[465];
	assign leaf[8316] = !f[743] && f[398] && f[344] && f[465];
	assign leaf[8317] = f[743] && !f[521];
	assign leaf[8318] = f[743] && f[521] && !f[411];
	assign leaf[8319] = f[743] && f[521] && f[411];
	
	// Tree 595, Classifier 5, Iteration: 59
	assign leaf[8320] = !f[442] && !f[538] && !f[160] && !f[546];
	assign leaf[8321] = !f[442] && !f[538] && !f[160] && f[546];
	assign leaf[8322] = !f[442] && !f[538] && f[160] && !f[513];
	assign leaf[8323] = !f[442] && !f[538] && f[160] && f[513];
	assign leaf[8324] = !f[442] && f[538] && !f[400] && !f[316];
	assign leaf[8325] = !f[442] && f[538] && !f[400] && f[316];
	assign leaf[8326] = !f[442] && f[538] && f[400] && !f[454];
	assign leaf[8327] = !f[442] && f[538] && f[400] && f[454];
	assign leaf[8328] = f[442] && !f[176] && !f[245] && !f[262];
	assign leaf[8329] = f[442] && !f[176] && !f[245] && f[262];
	assign leaf[8330] = f[442] && !f[176] && f[245] && !f[567];
	assign leaf[8331] = f[442] && !f[176] && f[245] && f[567];
	assign leaf[8332] = f[442] && f[176] && !f[179];
	assign leaf[8333] = f[442] && f[176] && f[179] && !f[287];
	assign leaf[8334] = f[442] && f[176] && f[179] && f[287];
	
	// Tree 596, Classifier 6, Iteration: 59
	assign leaf[8335] = !f[601] && !f[164] && !f[128] && !f[547];
	assign leaf[8336] = !f[601] && !f[164] && !f[128] && f[547];
	assign leaf[8337] = !f[601] && !f[164] && f[128] && !f[571];
	assign leaf[8338] = !f[601] && !f[164] && f[128] && f[571];
	assign leaf[8339] = !f[601] && f[164];
	assign leaf[8340] = f[601] && !f[129] && !f[238] && !f[627];
	assign leaf[8341] = f[601] && !f[129] && !f[238] && f[627];
	assign leaf[8342] = f[601] && !f[129] && f[238] && !f[99];
	assign leaf[8343] = f[601] && !f[129] && f[238] && f[99];
	assign leaf[8344] = f[601] && f[129] && !f[574] && !f[183];
	assign leaf[8345] = f[601] && f[129] && !f[574] && f[183];
	assign leaf[8346] = f[601] && f[129] && f[574] && !f[266];
	assign leaf[8347] = f[601] && f[129] && f[574] && f[266];
	
	// Tree 597, Classifier 7, Iteration: 59
	assign leaf[8348] = !f[129] && !f[122] && !f[432] && !f[377];
	assign leaf[8349] = !f[129] && !f[122] && !f[432] && f[377];
	assign leaf[8350] = !f[129] && !f[122] && f[432] && !f[345];
	assign leaf[8351] = !f[129] && !f[122] && f[432] && f[345];
	assign leaf[8352] = !f[129] && f[122];
	assign leaf[8353] = f[129];
	
	// Tree 598, Classifier 8, Iteration: 59
	assign leaf[8354] = !f[276] && !f[284] && !f[684] && !f[601];
	assign leaf[8355] = !f[276] && !f[284] && !f[684] && f[601];
	assign leaf[8356] = !f[276] && !f[284] && f[684] && !f[601];
	assign leaf[8357] = !f[276] && !f[284] && f[684] && f[601];
	assign leaf[8358] = !f[276] && f[284] && !f[374] && !f[354];
	assign leaf[8359] = !f[276] && f[284] && !f[374] && f[354];
	assign leaf[8360] = !f[276] && f[284] && f[374];
	assign leaf[8361] = f[276] && !f[403] && !f[543];
	assign leaf[8362] = f[276] && !f[403] && f[543] && !f[299];
	assign leaf[8363] = f[276] && !f[403] && f[543] && f[299];
	assign leaf[8364] = f[276] && f[403] && !f[207] && !f[511];
	assign leaf[8365] = f[276] && f[403] && !f[207] && f[511];
	assign leaf[8366] = f[276] && f[403] && f[207] && !f[682];
	assign leaf[8367] = f[276] && f[403] && f[207] && f[682];
	
	// Tree 599, Classifier 9, Iteration: 59
	assign leaf[8368] = !f[131] && !f[178] && !f[259] && !f[205];
	assign leaf[8369] = !f[131] && !f[178] && !f[259] && f[205];
	assign leaf[8370] = !f[131] && !f[178] && f[259] && !f[206];
	assign leaf[8371] = !f[131] && !f[178] && f[259] && f[206];
	assign leaf[8372] = !f[131] && f[178] && !f[181] && !f[691];
	assign leaf[8373] = !f[131] && f[178] && !f[181] && f[691];
	assign leaf[8374] = !f[131] && f[178] && f[181] && !f[210];
	assign leaf[8375] = !f[131] && f[178] && f[181] && f[210];
	assign leaf[8376] = f[131] && !f[128];
	assign leaf[8377] = f[131] && f[128];
	
	// Tree 600, Classifier 0, Iteration: 60
	assign leaf[8378] = !f[605] && !f[321] && !f[320] && !f[431];
	assign leaf[8379] = !f[605] && !f[321] && !f[320] && f[431];
	assign leaf[8380] = !f[605] && !f[321] && f[320] && !f[468];
	assign leaf[8381] = !f[605] && !f[321] && f[320] && f[468];
	assign leaf[8382] = !f[605] && f[321] && !f[153] && !f[480];
	assign leaf[8383] = !f[605] && f[321] && !f[153] && f[480];
	assign leaf[8384] = !f[605] && f[321] && f[153] && !f[401];
	assign leaf[8385] = !f[605] && f[321] && f[153] && f[401];
	assign leaf[8386] = f[605] && !f[207] && !f[492] && !f[273];
	assign leaf[8387] = f[605] && !f[207] && !f[492] && f[273];
	assign leaf[8388] = f[605] && !f[207] && f[492] && !f[128];
	assign leaf[8389] = f[605] && !f[207] && f[492] && f[128];
	assign leaf[8390] = f[605] && f[207] && !f[185] && !f[354];
	assign leaf[8391] = f[605] && f[207] && !f[185] && f[354];
	assign leaf[8392] = f[605] && f[207] && f[185] && !f[316];
	assign leaf[8393] = f[605] && f[207] && f[185] && f[316];
	
	// Tree 601, Classifier 1, Iteration: 60
	assign leaf[8394] = !f[710] && !f[716] && !f[181] && !f[125];
	assign leaf[8395] = !f[710] && !f[716] && !f[181] && f[125];
	assign leaf[8396] = !f[710] && !f[716] && f[181] && !f[266];
	assign leaf[8397] = !f[710] && !f[716] && f[181] && f[266];
	assign leaf[8398] = !f[710] && f[716];
	assign leaf[8399] = f[710];
	
	// Tree 602, Classifier 2, Iteration: 60
	assign leaf[8400] = !f[513] && !f[404] && !f[257] && !f[571];
	assign leaf[8401] = !f[513] && !f[404] && !f[257] && f[571];
	assign leaf[8402] = !f[513] && !f[404] && f[257] && !f[204];
	assign leaf[8403] = !f[513] && !f[404] && f[257] && f[204];
	assign leaf[8404] = !f[513] && f[404] && !f[483] && !f[241];
	assign leaf[8405] = !f[513] && f[404] && !f[483] && f[241];
	assign leaf[8406] = !f[513] && f[404] && f[483] && !f[401];
	assign leaf[8407] = !f[513] && f[404] && f[483] && f[401];
	assign leaf[8408] = f[513] && !f[433] && !f[381] && !f[454];
	assign leaf[8409] = f[513] && !f[433] && !f[381] && f[454];
	assign leaf[8410] = f[513] && !f[433] && f[381] && !f[295];
	assign leaf[8411] = f[513] && !f[433] && f[381] && f[295];
	assign leaf[8412] = f[513] && f[433] && !f[257] && !f[322];
	assign leaf[8413] = f[513] && f[433] && !f[257] && f[322];
	assign leaf[8414] = f[513] && f[433] && f[257] && !f[262];
	assign leaf[8415] = f[513] && f[433] && f[257] && f[262];
	
	// Tree 603, Classifier 3, Iteration: 60
	assign leaf[8416] = !f[429] && !f[127] && !f[209] && !f[173];
	assign leaf[8417] = !f[429] && !f[127] && !f[209] && f[173];
	assign leaf[8418] = !f[429] && !f[127] && f[209] && !f[320];
	assign leaf[8419] = !f[429] && !f[127] && f[209] && f[320];
	assign leaf[8420] = !f[429] && f[127] && !f[459] && !f[235];
	assign leaf[8421] = !f[429] && f[127] && !f[459] && f[235];
	assign leaf[8422] = !f[429] && f[127] && f[459] && !f[652];
	assign leaf[8423] = !f[429] && f[127] && f[459] && f[652];
	assign leaf[8424] = f[429] && !f[544] && !f[513] && !f[553];
	assign leaf[8425] = f[429] && !f[544] && !f[513] && f[553];
	assign leaf[8426] = f[429] && !f[544] && f[513] && !f[130];
	assign leaf[8427] = f[429] && !f[544] && f[513] && f[130];
	assign leaf[8428] = f[429] && f[544] && !f[687] && !f[549];
	assign leaf[8429] = f[429] && f[544] && !f[687] && f[549];
	assign leaf[8430] = f[429] && f[544] && f[687] && !f[327];
	assign leaf[8431] = f[429] && f[544] && f[687] && f[327];
	
	// Tree 604, Classifier 4, Iteration: 60
	assign leaf[8432] = !f[179] && !f[154] && !f[404] && !f[636];
	assign leaf[8433] = !f[179] && !f[154] && !f[404] && f[636];
	assign leaf[8434] = !f[179] && !f[154] && f[404] && !f[434];
	assign leaf[8435] = !f[179] && !f[154] && f[404] && f[434];
	assign leaf[8436] = !f[179] && f[154] && !f[156] && !f[128];
	assign leaf[8437] = !f[179] && f[154] && !f[156] && f[128];
	assign leaf[8438] = !f[179] && f[154] && f[156] && !f[266];
	assign leaf[8439] = !f[179] && f[154] && f[156] && f[266];
	assign leaf[8440] = f[179] && !f[235] && !f[405] && !f[180];
	assign leaf[8441] = f[179] && !f[235] && !f[405] && f[180];
	assign leaf[8442] = f[179] && !f[235] && f[405] && !f[262];
	assign leaf[8443] = f[179] && !f[235] && f[405] && f[262];
	assign leaf[8444] = f[179] && f[235] && !f[214] && !f[181];
	assign leaf[8445] = f[179] && f[235] && !f[214] && f[181];
	assign leaf[8446] = f[179] && f[235] && f[214] && !f[155];
	assign leaf[8447] = f[179] && f[235] && f[214] && f[155];
	
	// Tree 605, Classifier 5, Iteration: 60
	assign leaf[8448] = !f[713] && !f[630] && !f[403] && !f[511];
	assign leaf[8449] = !f[713] && !f[630] && !f[403] && f[511];
	assign leaf[8450] = !f[713] && !f[630] && f[403] && !f[406];
	assign leaf[8451] = !f[713] && !f[630] && f[403] && f[406];
	assign leaf[8452] = !f[713] && f[630] && !f[347] && !f[270];
	assign leaf[8453] = !f[713] && f[630] && !f[347] && f[270];
	assign leaf[8454] = !f[713] && f[630] && f[347] && !f[263];
	assign leaf[8455] = !f[713] && f[630] && f[347] && f[263];
	assign leaf[8456] = f[713] && !f[574] && !f[240] && !f[460];
	assign leaf[8457] = f[713] && !f[574] && !f[240] && f[460];
	assign leaf[8458] = f[713] && !f[574] && f[240] && !f[434];
	assign leaf[8459] = f[713] && !f[574] && f[240] && f[434];
	assign leaf[8460] = f[713] && f[574] && !f[710] && !f[683];
	assign leaf[8461] = f[713] && f[574] && !f[710] && f[683];
	assign leaf[8462] = f[713] && f[574] && f[710];
	
	// Tree 606, Classifier 6, Iteration: 60
	assign leaf[8463] = !f[205] && !f[467] && !f[326] && !f[123];
	assign leaf[8464] = !f[205] && !f[467] && !f[326] && f[123];
	assign leaf[8465] = !f[205] && !f[467] && f[326] && !f[469];
	assign leaf[8466] = !f[205] && !f[467] && f[326] && f[469];
	assign leaf[8467] = !f[205] && f[467] && !f[432] && !f[436];
	assign leaf[8468] = !f[205] && f[467] && !f[432] && f[436];
	assign leaf[8469] = !f[205] && f[467] && f[432] && !f[287];
	assign leaf[8470] = !f[205] && f[467] && f[432] && f[287];
	assign leaf[8471] = f[205] && !f[348] && !f[183] && !f[294];
	assign leaf[8472] = f[205] && !f[348] && !f[183] && f[294];
	assign leaf[8473] = f[205] && !f[348] && f[183] && !f[573];
	assign leaf[8474] = f[205] && !f[348] && f[183] && f[573];
	assign leaf[8475] = f[205] && f[348] && !f[344] && !f[325];
	assign leaf[8476] = f[205] && f[348] && !f[344] && f[325];
	assign leaf[8477] = f[205] && f[348] && f[344] && !f[488];
	assign leaf[8478] = f[205] && f[348] && f[344] && f[488];
	
	// Tree 607, Classifier 7, Iteration: 60
	assign leaf[8479] = !f[239] && !f[236] && !f[327] && !f[156];
	assign leaf[8480] = !f[239] && !f[236] && !f[327] && f[156];
	assign leaf[8481] = !f[239] && !f[236] && f[327] && !f[206];
	assign leaf[8482] = !f[239] && !f[236] && f[327] && f[206];
	assign leaf[8483] = !f[239] && f[236] && !f[247] && !f[685];
	assign leaf[8484] = !f[239] && f[236] && !f[247] && f[685];
	assign leaf[8485] = !f[239] && f[236] && f[247];
	assign leaf[8486] = f[239] && !f[371] && !f[369] && !f[457];
	assign leaf[8487] = f[239] && !f[371] && !f[369] && f[457];
	assign leaf[8488] = f[239] && !f[371] && f[369] && !f[489];
	assign leaf[8489] = f[239] && !f[371] && f[369] && f[489];
	assign leaf[8490] = f[239] && f[371] && !f[460] && !f[293];
	assign leaf[8491] = f[239] && f[371] && !f[460] && f[293];
	assign leaf[8492] = f[239] && f[371] && f[460] && !f[428];
	assign leaf[8493] = f[239] && f[371] && f[460] && f[428];
	
	// Tree 608, Classifier 8, Iteration: 60
	assign leaf[8494] = !f[469] && !f[317] && !f[627] && !f[653];
	assign leaf[8495] = !f[469] && !f[317] && !f[627] && f[653];
	assign leaf[8496] = !f[469] && !f[317] && f[627] && !f[600];
	assign leaf[8497] = !f[469] && !f[317] && f[627] && f[600];
	assign leaf[8498] = !f[469] && f[317] && !f[375] && !f[430];
	assign leaf[8499] = !f[469] && f[317] && !f[375] && f[430];
	assign leaf[8500] = !f[469] && f[317] && f[375] && !f[401];
	assign leaf[8501] = !f[469] && f[317] && f[375] && f[401];
	assign leaf[8502] = f[469] && !f[523] && !f[180] && !f[569];
	assign leaf[8503] = f[469] && !f[523] && !f[180] && f[569];
	assign leaf[8504] = f[469] && !f[523] && f[180] && !f[314];
	assign leaf[8505] = f[469] && !f[523] && f[180] && f[314];
	assign leaf[8506] = f[469] && f[523] && !f[218] && !f[638];
	assign leaf[8507] = f[469] && f[523] && !f[218] && f[638];
	assign leaf[8508] = f[469] && f[523] && f[218] && !f[574];
	assign leaf[8509] = f[469] && f[523] && f[218] && f[574];
	
	// Tree 609, Classifier 9, Iteration: 60
	assign leaf[8510] = !f[709] && !f[627] && !f[404] && !f[182];
	assign leaf[8511] = !f[709] && !f[627] && !f[404] && f[182];
	assign leaf[8512] = !f[709] && !f[627] && f[404] && !f[378];
	assign leaf[8513] = !f[709] && !f[627] && f[404] && f[378];
	assign leaf[8514] = !f[709] && f[627] && !f[516] && !f[485];
	assign leaf[8515] = !f[709] && f[627] && !f[516] && f[485];
	assign leaf[8516] = !f[709] && f[627] && f[516] && !f[186];
	assign leaf[8517] = !f[709] && f[627] && f[516] && f[186];
	assign leaf[8518] = f[709] && !f[264] && !f[293] && !f[316];
	assign leaf[8519] = f[709] && !f[264] && !f[293] && f[316];
	assign leaf[8520] = f[709] && !f[264] && f[293] && !f[375];
	assign leaf[8521] = f[709] && !f[264] && f[293] && f[375];
	assign leaf[8522] = f[709] && f[264] && !f[213] && !f[268];
	assign leaf[8523] = f[709] && f[264] && !f[213] && f[268];
	assign leaf[8524] = f[709] && f[264] && f[213] && !f[712];
	assign leaf[8525] = f[709] && f[264] && f[213] && f[712];
	
	// Tree 610, Classifier 0, Iteration: 61
	assign leaf[8526] = !f[572] && !f[547] && !f[376] && !f[460];
	assign leaf[8527] = !f[572] && !f[547] && !f[376] && f[460];
	assign leaf[8528] = !f[572] && !f[547] && f[376] && !f[189];
	assign leaf[8529] = !f[572] && !f[547] && f[376] && f[189];
	assign leaf[8530] = !f[572] && f[547] && !f[294] && !f[268];
	assign leaf[8531] = !f[572] && f[547] && !f[294] && f[268];
	assign leaf[8532] = !f[572] && f[547] && f[294] && !f[576];
	assign leaf[8533] = !f[572] && f[547] && f[294] && f[576];
	assign leaf[8534] = f[572] && !f[683] && !f[319] && !f[354];
	assign leaf[8535] = f[572] && !f[683] && !f[319] && f[354];
	assign leaf[8536] = f[572] && !f[683] && f[319] && !f[598];
	assign leaf[8537] = f[572] && !f[683] && f[319] && f[598];
	assign leaf[8538] = f[572] && f[683];
	
	// Tree 611, Classifier 1, Iteration: 61
	assign leaf[8539] = !f[204] && !f[634] && !f[493] && !f[235];
	assign leaf[8540] = !f[204] && !f[634] && !f[493] && f[235];
	assign leaf[8541] = !f[204] && !f[634] && f[493] && !f[547];
	assign leaf[8542] = !f[204] && !f[634] && f[493] && f[547];
	assign leaf[8543] = !f[204] && f[634] && !f[348] && !f[654];
	assign leaf[8544] = !f[204] && f[634] && !f[348] && f[654];
	assign leaf[8545] = !f[204] && f[634] && f[348] && !f[157];
	assign leaf[8546] = !f[204] && f[634] && f[348] && f[157];
	assign leaf[8547] = f[204] && !f[544] && !f[599] && !f[575];
	assign leaf[8548] = f[204] && !f[544] && !f[599] && f[575];
	assign leaf[8549] = f[204] && !f[544] && f[599];
	assign leaf[8550] = f[204] && f[544] && !f[609];
	assign leaf[8551] = f[204] && f[544] && f[609];
	
	// Tree 612, Classifier 2, Iteration: 61
	assign leaf[8552] = !f[351] && !f[547] && !f[261] && !f[681];
	assign leaf[8553] = !f[351] && !f[547] && !f[261] && f[681];
	assign leaf[8554] = !f[351] && !f[547] && f[261] && !f[657];
	assign leaf[8555] = !f[351] && !f[547] && f[261] && f[657];
	assign leaf[8556] = !f[351] && f[547] && !f[407] && !f[512];
	assign leaf[8557] = !f[351] && f[547] && !f[407] && f[512];
	assign leaf[8558] = !f[351] && f[547] && f[407] && !f[630];
	assign leaf[8559] = !f[351] && f[547] && f[407] && f[630];
	assign leaf[8560] = f[351] && !f[437] && !f[605] && !f[524];
	assign leaf[8561] = f[351] && !f[437] && !f[605] && f[524];
	assign leaf[8562] = f[351] && !f[437] && f[605] && !f[520];
	assign leaf[8563] = f[351] && !f[437] && f[605] && f[520];
	assign leaf[8564] = f[351] && f[437] && !f[659] && !f[482];
	assign leaf[8565] = f[351] && f[437] && !f[659] && f[482];
	assign leaf[8566] = f[351] && f[437] && f[659] && !f[257];
	assign leaf[8567] = f[351] && f[437] && f[659] && f[257];
	
	// Tree 613, Classifier 3, Iteration: 61
	assign leaf[8568] = !f[384] && !f[358] && !f[328] && !f[190];
	assign leaf[8569] = !f[384] && !f[358] && !f[328] && f[190];
	assign leaf[8570] = !f[384] && !f[358] && f[328] && !f[241];
	assign leaf[8571] = !f[384] && !f[358] && f[328] && f[241];
	assign leaf[8572] = !f[384] && f[358];
	assign leaf[8573] = f[384] && !f[266] && !f[131] && !f[461];
	assign leaf[8574] = f[384] && !f[266] && !f[131] && f[461];
	assign leaf[8575] = f[384] && !f[266] && f[131] && !f[236];
	assign leaf[8576] = f[384] && !f[266] && f[131] && f[236];
	assign leaf[8577] = f[384] && f[266] && !f[122] && !f[298];
	assign leaf[8578] = f[384] && f[266] && !f[122] && f[298];
	assign leaf[8579] = f[384] && f[266] && f[122] && !f[261];
	assign leaf[8580] = f[384] && f[266] && f[122] && f[261];
	
	// Tree 614, Classifier 4, Iteration: 61
	assign leaf[8581] = !f[519] && !f[630] && !f[686] && !f[201];
	assign leaf[8582] = !f[519] && !f[630] && !f[686] && f[201];
	assign leaf[8583] = !f[519] && !f[630] && f[686] && !f[660];
	assign leaf[8584] = !f[519] && !f[630] && f[686] && f[660];
	assign leaf[8585] = !f[519] && f[630] && !f[605] && !f[181];
	assign leaf[8586] = !f[519] && f[630] && !f[605] && f[181];
	assign leaf[8587] = !f[519] && f[630] && f[605] && !f[328];
	assign leaf[8588] = !f[519] && f[630] && f[605] && f[328];
	assign leaf[8589] = f[519] && !f[524] && !f[186] && !f[297];
	assign leaf[8590] = f[519] && !f[524] && !f[186] && f[297];
	assign leaf[8591] = f[519] && !f[524] && f[186] && !f[269];
	assign leaf[8592] = f[519] && !f[524] && f[186] && f[269];
	assign leaf[8593] = f[519] && f[524] && !f[261] && !f[387];
	assign leaf[8594] = f[519] && f[524] && !f[261] && f[387];
	assign leaf[8595] = f[519] && f[524] && f[261] && !f[273];
	assign leaf[8596] = f[519] && f[524] && f[261] && f[273];
	
	// Tree 615, Classifier 5, Iteration: 61
	assign leaf[8597] = !f[459] && !f[411] && !f[551] && !f[151];
	assign leaf[8598] = !f[459] && !f[411] && !f[551] && f[151];
	assign leaf[8599] = !f[459] && !f[411] && f[551] && !f[294];
	assign leaf[8600] = !f[459] && !f[411] && f[551] && f[294];
	assign leaf[8601] = !f[459] && f[411] && !f[329] && !f[179];
	assign leaf[8602] = !f[459] && f[411] && !f[329] && f[179];
	assign leaf[8603] = !f[459] && f[411] && f[329];
	assign leaf[8604] = f[459] && !f[430] && !f[712] && !f[375];
	assign leaf[8605] = f[459] && !f[430] && !f[712] && f[375];
	assign leaf[8606] = f[459] && !f[430] && f[712];
	assign leaf[8607] = f[459] && f[430] && !f[542] && !f[627];
	assign leaf[8608] = f[459] && f[430] && !f[542] && f[627];
	assign leaf[8609] = f[459] && f[430] && f[542] && !f[576];
	assign leaf[8610] = f[459] && f[430] && f[542] && f[576];
	
	// Tree 616, Classifier 6, Iteration: 61
	assign leaf[8611] = !f[541] && !f[516] && !f[511] && !f[514];
	assign leaf[8612] = !f[541] && !f[516] && !f[511] && f[514];
	assign leaf[8613] = !f[541] && !f[516] && f[511] && !f[600];
	assign leaf[8614] = !f[541] && !f[516] && f[511] && f[600];
	assign leaf[8615] = !f[541] && f[516] && !f[575] && !f[571];
	assign leaf[8616] = !f[541] && f[516] && !f[575] && f[571];
	assign leaf[8617] = !f[541] && f[516] && f[575] && !f[485];
	assign leaf[8618] = !f[541] && f[516] && f[575] && f[485];
	assign leaf[8619] = f[541] && !f[401] && !f[291] && !f[237];
	assign leaf[8620] = f[541] && !f[401] && !f[291] && f[237];
	assign leaf[8621] = f[541] && !f[401] && f[291] && !f[371];
	assign leaf[8622] = f[541] && !f[401] && f[291] && f[371];
	assign leaf[8623] = f[541] && f[401] && !f[457] && !f[403];
	assign leaf[8624] = f[541] && f[401] && !f[457] && f[403];
	assign leaf[8625] = f[541] && f[401] && f[457] && !f[136];
	assign leaf[8626] = f[541] && f[401] && f[457] && f[136];
	
	// Tree 617, Classifier 7, Iteration: 61
	assign leaf[8627] = !f[582] && !f[161] && !f[272] && !f[355];
	assign leaf[8628] = !f[582] && !f[161] && !f[272] && f[355];
	assign leaf[8629] = !f[582] && !f[161] && f[272] && !f[406];
	assign leaf[8630] = !f[582] && !f[161] && f[272] && f[406];
	assign leaf[8631] = !f[582] && f[161];
	assign leaf[8632] = f[582] && !f[350] && !f[212];
	assign leaf[8633] = f[582] && !f[350] && f[212];
	assign leaf[8634] = f[582] && f[350];
	
	// Tree 618, Classifier 8, Iteration: 61
	assign leaf[8635] = !f[466] && !f[549] && !f[575] && !f[324];
	assign leaf[8636] = !f[466] && !f[549] && !f[575] && f[324];
	assign leaf[8637] = !f[466] && !f[549] && f[575] && !f[659];
	assign leaf[8638] = !f[466] && !f[549] && f[575] && f[659];
	assign leaf[8639] = !f[466] && f[549] && !f[576] && !f[523];
	assign leaf[8640] = !f[466] && f[549] && !f[576] && f[523];
	assign leaf[8641] = !f[466] && f[549] && f[576] && !f[178];
	assign leaf[8642] = !f[466] && f[549] && f[576] && f[178];
	assign leaf[8643] = f[466] && !f[520] && !f[436] && !f[267];
	assign leaf[8644] = f[466] && !f[520] && !f[436] && f[267];
	assign leaf[8645] = f[466] && !f[520] && f[436] && !f[351];
	assign leaf[8646] = f[466] && !f[520] && f[436] && f[351];
	assign leaf[8647] = f[466] && f[520] && !f[284] && !f[594];
	assign leaf[8648] = f[466] && f[520] && !f[284] && f[594];
	assign leaf[8649] = f[466] && f[520] && f[284];
	
	// Tree 619, Classifier 9, Iteration: 61
	assign leaf[8650] = !f[740] && !f[462] && !f[457] && !f[181];
	assign leaf[8651] = !f[740] && !f[462] && !f[457] && f[181];
	assign leaf[8652] = !f[740] && !f[462] && f[457] && !f[375];
	assign leaf[8653] = !f[740] && !f[462] && f[457] && f[375];
	assign leaf[8654] = !f[740] && f[462] && !f[401] && !f[427];
	assign leaf[8655] = !f[740] && f[462] && !f[401] && f[427];
	assign leaf[8656] = !f[740] && f[462] && f[401] && !f[290];
	assign leaf[8657] = !f[740] && f[462] && f[401] && f[290];
	assign leaf[8658] = f[740] && !f[240] && !f[272];
	assign leaf[8659] = f[740] && !f[240] && f[272];
	assign leaf[8660] = f[740] && f[240] && !f[214] && !f[437];
	assign leaf[8661] = f[740] && f[240] && !f[214] && f[437];
	assign leaf[8662] = f[740] && f[240] && f[214] && !f[410];
	assign leaf[8663] = f[740] && f[240] && f[214] && f[410];
	
	// Tree 620, Classifier 0, Iteration: 62
	assign leaf[8664] = !f[572] && !f[541] && !f[494] && !f[595];
	assign leaf[8665] = !f[572] && !f[541] && !f[494] && f[595];
	assign leaf[8666] = !f[572] && !f[541] && f[494] && !f[316];
	assign leaf[8667] = !f[572] && !f[541] && f[494] && f[316];
	assign leaf[8668] = !f[572] && f[541] && !f[353] && !f[485];
	assign leaf[8669] = !f[572] && f[541] && !f[353] && f[485];
	assign leaf[8670] = !f[572] && f[541] && f[353] && !f[607];
	assign leaf[8671] = !f[572] && f[541] && f[353] && f[607];
	assign leaf[8672] = f[572] && !f[683] && !f[459] && !f[455];
	assign leaf[8673] = f[572] && !f[683] && !f[459] && f[455];
	assign leaf[8674] = f[572] && !f[683] && f[459] && !f[686];
	assign leaf[8675] = f[572] && !f[683] && f[459] && f[686];
	assign leaf[8676] = f[572] && f[683] && !f[549];
	assign leaf[8677] = f[572] && f[683] && f[549];
	
	// Tree 621, Classifier 1, Iteration: 62
	assign leaf[8678] = !f[381] && !f[242] && !f[155] && !f[295];
	assign leaf[8679] = !f[381] && !f[242] && !f[155] && f[295];
	assign leaf[8680] = !f[381] && !f[242] && f[155] && !f[465];
	assign leaf[8681] = !f[381] && !f[242] && f[155] && f[465];
	assign leaf[8682] = !f[381] && f[242] && !f[519] && !f[183];
	assign leaf[8683] = !f[381] && f[242] && !f[519] && f[183];
	assign leaf[8684] = !f[381] && f[242] && f[519] && !f[408];
	assign leaf[8685] = !f[381] && f[242] && f[519] && f[408];
	assign leaf[8686] = f[381] && !f[297] && !f[576] && !f[460];
	assign leaf[8687] = f[381] && !f[297] && !f[576] && f[460];
	assign leaf[8688] = f[381] && !f[297] && f[576] && !f[125];
	assign leaf[8689] = f[381] && !f[297] && f[576] && f[125];
	assign leaf[8690] = f[381] && f[297] && !f[463] && !f[238];
	assign leaf[8691] = f[381] && f[297] && !f[463] && f[238];
	assign leaf[8692] = f[381] && f[297] && f[463] && !f[207];
	assign leaf[8693] = f[381] && f[297] && f[463] && f[207];
	
	// Tree 622, Classifier 2, Iteration: 62
	assign leaf[8694] = !f[121] && !f[497] && !f[607] && !f[689];
	assign leaf[8695] = !f[121] && !f[497] && !f[607] && f[689];
	assign leaf[8696] = !f[121] && !f[497] && f[607] && !f[551];
	assign leaf[8697] = !f[121] && !f[497] && f[607] && f[551];
	assign leaf[8698] = !f[121] && f[497] && !f[633] && !f[609];
	assign leaf[8699] = !f[121] && f[497] && !f[633] && f[609];
	assign leaf[8700] = !f[121] && f[497] && f[633] && !f[353];
	assign leaf[8701] = !f[121] && f[497] && f[633] && f[353];
	assign leaf[8702] = f[121] && !f[232] && !f[605];
	assign leaf[8703] = f[121] && !f[232] && f[605] && !f[608];
	assign leaf[8704] = f[121] && !f[232] && f[605] && f[608];
	assign leaf[8705] = f[121] && f[232] && !f[467];
	assign leaf[8706] = f[121] && f[232] && f[467];
	
	// Tree 623, Classifier 3, Iteration: 62
	assign leaf[8707] = !f[705] && !f[386] && !f[346] && !f[372];
	assign leaf[8708] = !f[705] && !f[386] && !f[346] && f[372];
	assign leaf[8709] = !f[705] && !f[386] && f[346] && !f[321];
	assign leaf[8710] = !f[705] && !f[386] && f[346] && f[321];
	assign leaf[8711] = !f[705] && f[386] && !f[152] && !f[508];
	assign leaf[8712] = !f[705] && f[386] && !f[152] && f[508];
	assign leaf[8713] = !f[705] && f[386] && f[152] && !f[237];
	assign leaf[8714] = !f[705] && f[386] && f[152] && f[237];
	assign leaf[8715] = f[705];
	
	// Tree 624, Classifier 4, Iteration: 62
	assign leaf[8716] = !f[318] && !f[320] && !f[316] && !f[257];
	assign leaf[8717] = !f[318] && !f[320] && !f[316] && f[257];
	assign leaf[8718] = !f[318] && !f[320] && f[316] && !f[264];
	assign leaf[8719] = !f[318] && !f[320] && f[316] && f[264];
	assign leaf[8720] = !f[318] && f[320] && !f[262] && !f[274];
	assign leaf[8721] = !f[318] && f[320] && !f[262] && f[274];
	assign leaf[8722] = !f[318] && f[320] && f[262] && !f[577];
	assign leaf[8723] = !f[318] && f[320] && f[262] && f[577];
	assign leaf[8724] = f[318] && !f[321] && !f[237] && !f[181];
	assign leaf[8725] = f[318] && !f[321] && !f[237] && f[181];
	assign leaf[8726] = f[318] && !f[321] && f[237] && !f[320];
	assign leaf[8727] = f[318] && !f[321] && f[237] && f[320];
	assign leaf[8728] = f[318] && f[321] && !f[183] && !f[289];
	assign leaf[8729] = f[318] && f[321] && !f[183] && f[289];
	assign leaf[8730] = f[318] && f[321] && f[183] && !f[296];
	assign leaf[8731] = f[318] && f[321] && f[183] && f[296];
	
	// Tree 625, Classifier 5, Iteration: 62
	assign leaf[8732] = !f[402] && !f[630] && !f[270] && !f[126];
	assign leaf[8733] = !f[402] && !f[630] && !f[270] && f[126];
	assign leaf[8734] = !f[402] && !f[630] && f[270] && !f[214];
	assign leaf[8735] = !f[402] && !f[630] && f[270] && f[214];
	assign leaf[8736] = !f[402] && f[630] && !f[269] && !f[157];
	assign leaf[8737] = !f[402] && f[630] && !f[269] && f[157];
	assign leaf[8738] = !f[402] && f[630] && f[269] && !f[265];
	assign leaf[8739] = !f[402] && f[630] && f[269] && f[265];
	assign leaf[8740] = f[402] && !f[546] && !f[344] && !f[294];
	assign leaf[8741] = f[402] && !f[546] && !f[344] && f[294];
	assign leaf[8742] = f[402] && !f[546] && f[344] && !f[427];
	assign leaf[8743] = f[402] && !f[546] && f[344] && f[427];
	assign leaf[8744] = f[402] && f[546] && !f[185] && !f[234];
	assign leaf[8745] = f[402] && f[546] && !f[185] && f[234];
	assign leaf[8746] = f[402] && f[546] && f[185] && !f[378];
	assign leaf[8747] = f[402] && f[546] && f[185] && f[378];
	
	// Tree 626, Classifier 6, Iteration: 62
	assign leaf[8748] = !f[297] && !f[656] && !f[217] && !f[350];
	assign leaf[8749] = !f[297] && !f[656] && !f[217] && f[350];
	assign leaf[8750] = !f[297] && !f[656] && f[217] && !f[580];
	assign leaf[8751] = !f[297] && !f[656] && f[217] && f[580];
	assign leaf[8752] = !f[297] && f[656] && !f[355] && !f[152];
	assign leaf[8753] = !f[297] && f[656] && !f[355] && f[152];
	assign leaf[8754] = !f[297] && f[656] && f[355] && !f[125];
	assign leaf[8755] = !f[297] && f[656] && f[355] && f[125];
	assign leaf[8756] = f[297] && !f[573] && !f[359] && !f[287];
	assign leaf[8757] = f[297] && !f[573] && !f[359] && f[287];
	assign leaf[8758] = f[297] && !f[573] && f[359];
	assign leaf[8759] = f[297] && f[573] && !f[350] && !f[273];
	assign leaf[8760] = f[297] && f[573] && !f[350] && f[273];
	assign leaf[8761] = f[297] && f[573] && f[350] && !f[212];
	assign leaf[8762] = f[297] && f[573] && f[350] && f[212];
	
	// Tree 627, Classifier 7, Iteration: 62
	assign leaf[8763] = !f[638] && !f[348] && !f[374] && !f[185];
	assign leaf[8764] = !f[638] && !f[348] && !f[374] && f[185];
	assign leaf[8765] = !f[638] && !f[348] && f[374] && !f[460];
	assign leaf[8766] = !f[638] && !f[348] && f[374] && f[460];
	assign leaf[8767] = !f[638] && f[348] && !f[401] && !f[210];
	assign leaf[8768] = !f[638] && f[348] && !f[401] && f[210];
	assign leaf[8769] = !f[638] && f[348] && f[401] && !f[460];
	assign leaf[8770] = !f[638] && f[348] && f[401] && f[460];
	assign leaf[8771] = f[638];
	
	// Tree 628, Classifier 8, Iteration: 62
	assign leaf[8772] = !f[437] && !f[291] && !f[657] && !f[573];
	assign leaf[8773] = !f[437] && !f[291] && !f[657] && f[573];
	assign leaf[8774] = !f[437] && !f[291] && f[657] && !f[517];
	assign leaf[8775] = !f[437] && !f[291] && f[657] && f[517];
	assign leaf[8776] = !f[437] && f[291] && !f[520] && !f[300];
	assign leaf[8777] = !f[437] && f[291] && !f[520] && f[300];
	assign leaf[8778] = !f[437] && f[291] && f[520] && !f[351];
	assign leaf[8779] = !f[437] && f[291] && f[520] && f[351];
	assign leaf[8780] = f[437] && !f[381] && !f[494] && !f[406];
	assign leaf[8781] = f[437] && !f[381] && !f[494] && f[406];
	assign leaf[8782] = f[437] && !f[381] && f[494] && !f[351];
	assign leaf[8783] = f[437] && !f[381] && f[494] && f[351];
	assign leaf[8784] = f[437] && f[381] && !f[273] && !f[179];
	assign leaf[8785] = f[437] && f[381] && !f[273] && f[179];
	assign leaf[8786] = f[437] && f[381] && f[273] && !f[686];
	assign leaf[8787] = f[437] && f[381] && f[273] && f[686];
	
	// Tree 629, Classifier 9, Iteration: 62
	assign leaf[8788] = !f[350] && !f[717] && !f[719] && !f[606];
	assign leaf[8789] = !f[350] && !f[717] && !f[719] && f[606];
	assign leaf[8790] = !f[350] && !f[717] && f[719] && !f[461];
	assign leaf[8791] = !f[350] && !f[717] && f[719] && f[461];
	assign leaf[8792] = !f[350] && f[717] && !f[237] && !f[608];
	assign leaf[8793] = !f[350] && f[717] && !f[237] && f[608];
	assign leaf[8794] = !f[350] && f[717] && f[237] && !f[378];
	assign leaf[8795] = !f[350] && f[717] && f[237] && f[378];
	assign leaf[8796] = f[350] && !f[488] && !f[324] && !f[373];
	assign leaf[8797] = f[350] && !f[488] && !f[324] && f[373];
	assign leaf[8798] = f[350] && !f[488] && f[324] && !f[187];
	assign leaf[8799] = f[350] && !f[488] && f[324] && f[187];
	assign leaf[8800] = f[350] && f[488] && !f[708] && !f[610];
	assign leaf[8801] = f[350] && f[488] && !f[708] && f[610];
	assign leaf[8802] = f[350] && f[488] && f[708] && !f[405];
	assign leaf[8803] = f[350] && f[488] && f[708] && f[405];
	
	// Tree 630, Classifier 0, Iteration: 63
	assign leaf[8804] = !f[380] && !f[382] && !f[303] && !f[517];
	assign leaf[8805] = !f[380] && !f[382] && !f[303] && f[517];
	assign leaf[8806] = !f[380] && !f[382] && f[303] && !f[385];
	assign leaf[8807] = !f[380] && !f[382] && f[303] && f[385];
	assign leaf[8808] = !f[380] && f[382] && !f[403] && !f[385];
	assign leaf[8809] = !f[380] && f[382] && !f[403] && f[385];
	assign leaf[8810] = !f[380] && f[382] && f[403] && !f[408];
	assign leaf[8811] = !f[380] && f[382] && f[403] && f[408];
	assign leaf[8812] = f[380] && !f[406] && !f[656] && !f[155];
	assign leaf[8813] = f[380] && !f[406] && !f[656] && f[155];
	assign leaf[8814] = f[380] && !f[406] && f[656] && !f[492];
	assign leaf[8815] = f[380] && !f[406] && f[656] && f[492];
	assign leaf[8816] = f[380] && f[406] && !f[244];
	assign leaf[8817] = f[380] && f[406] && f[244] && !f[129];
	assign leaf[8818] = f[380] && f[406] && f[244] && f[129];
	
	// Tree 631, Classifier 1, Iteration: 63
	assign leaf[8819] = !f[510] && !f[538] && !f[408] && !f[520];
	assign leaf[8820] = !f[510] && !f[538] && !f[408] && f[520];
	assign leaf[8821] = !f[510] && !f[538] && f[408] && !f[491];
	assign leaf[8822] = !f[510] && !f[538] && f[408] && f[491];
	assign leaf[8823] = !f[510] && f[538] && !f[625];
	assign leaf[8824] = !f[510] && f[538] && f[625];
	assign leaf[8825] = f[510];
	
	// Tree 632, Classifier 2, Iteration: 63
	assign leaf[8826] = !f[709] && !f[409] && !f[460] && !f[494];
	assign leaf[8827] = !f[709] && !f[409] && !f[460] && f[494];
	assign leaf[8828] = !f[709] && !f[409] && f[460] && !f[374];
	assign leaf[8829] = !f[709] && !f[409] && f[460] && f[374];
	assign leaf[8830] = !f[709] && f[409] && !f[463] && !f[491];
	assign leaf[8831] = !f[709] && f[409] && !f[463] && f[491];
	assign leaf[8832] = !f[709] && f[409] && f[463] && !f[679];
	assign leaf[8833] = !f[709] && f[409] && f[463] && f[679];
	assign leaf[8834] = f[709];
	
	// Tree 633, Classifier 3, Iteration: 63
	assign leaf[8835] = !f[707] && !f[571] && !f[546] && !f[490];
	assign leaf[8836] = !f[707] && !f[571] && !f[546] && f[490];
	assign leaf[8837] = !f[707] && !f[571] && f[546] && !f[492];
	assign leaf[8838] = !f[707] && !f[571] && f[546] && f[492];
	assign leaf[8839] = !f[707] && f[571] && !f[596] && !f[580];
	assign leaf[8840] = !f[707] && f[571] && !f[596] && f[580];
	assign leaf[8841] = !f[707] && f[571] && f[596] && !f[519];
	assign leaf[8842] = !f[707] && f[571] && f[596] && f[519];
	assign leaf[8843] = f[707] && !f[267];
	assign leaf[8844] = f[707] && f[267] && !f[571];
	assign leaf[8845] = f[707] && f[267] && f[571];
	
	// Tree 634, Classifier 4, Iteration: 63
	assign leaf[8846] = !f[381] && !f[515] && !f[321] && !f[182];
	assign leaf[8847] = !f[381] && !f[515] && !f[321] && f[182];
	assign leaf[8848] = !f[381] && !f[515] && f[321] && !f[662];
	assign leaf[8849] = !f[381] && !f[515] && f[321] && f[662];
	assign leaf[8850] = !f[381] && f[515] && !f[409] && !f[579];
	assign leaf[8851] = !f[381] && f[515] && !f[409] && f[579];
	assign leaf[8852] = !f[381] && f[515] && f[409] && !f[154];
	assign leaf[8853] = !f[381] && f[515] && f[409] && f[154];
	assign leaf[8854] = f[381] && !f[465] && !f[158] && !f[466];
	assign leaf[8855] = f[381] && !f[465] && !f[158] && f[466];
	assign leaf[8856] = f[381] && !f[465] && f[158] && !f[372];
	assign leaf[8857] = f[381] && !f[465] && f[158] && f[372];
	assign leaf[8858] = f[381] && f[465] && !f[235] && !f[316];
	assign leaf[8859] = f[381] && f[465] && !f[235] && f[316];
	assign leaf[8860] = f[381] && f[465] && f[235] && !f[246];
	assign leaf[8861] = f[381] && f[465] && f[235] && f[246];
	
	// Tree 635, Classifier 5, Iteration: 63
	assign leaf[8862] = !f[631] && !f[715] && !f[514] && !f[440];
	assign leaf[8863] = !f[631] && !f[715] && !f[514] && f[440];
	assign leaf[8864] = !f[631] && !f[715] && f[514] && !f[655];
	assign leaf[8865] = !f[631] && !f[715] && f[514] && f[655];
	assign leaf[8866] = !f[631] && f[715] && !f[463] && !f[294];
	assign leaf[8867] = !f[631] && f[715] && !f[463] && f[294];
	assign leaf[8868] = !f[631] && f[715] && f[463];
	assign leaf[8869] = f[631] && !f[457] && !f[159] && !f[553];
	assign leaf[8870] = f[631] && !f[457] && !f[159] && f[553];
	assign leaf[8871] = f[631] && !f[457] && f[159] && !f[211];
	assign leaf[8872] = f[631] && !f[457] && f[159] && f[211];
	assign leaf[8873] = f[631] && f[457] && !f[712] && !f[398];
	assign leaf[8874] = f[631] && f[457] && !f[712] && f[398];
	assign leaf[8875] = f[631] && f[457] && f[712] && !f[295];
	assign leaf[8876] = f[631] && f[457] && f[712] && f[295];
	
	// Tree 636, Classifier 6, Iteration: 63
	assign leaf[8877] = !f[268] && !f[349] && !f[686] && !f[322];
	assign leaf[8878] = !f[268] && !f[349] && !f[686] && f[322];
	assign leaf[8879] = !f[268] && !f[349] && f[686] && !f[546];
	assign leaf[8880] = !f[268] && !f[349] && f[686] && f[546];
	assign leaf[8881] = !f[268] && f[349] && !f[123] && !f[629];
	assign leaf[8882] = !f[268] && f[349] && !f[123] && f[629];
	assign leaf[8883] = !f[268] && f[349] && f[123] && !f[599];
	assign leaf[8884] = !f[268] && f[349] && f[123] && f[599];
	assign leaf[8885] = f[268] && !f[408] && !f[570] && !f[239];
	assign leaf[8886] = f[268] && !f[408] && !f[570] && f[239];
	assign leaf[8887] = f[268] && !f[408] && f[570] && !f[490];
	assign leaf[8888] = f[268] && !f[408] && f[570] && f[490];
	assign leaf[8889] = f[268] && f[408] && !f[349] && !f[606];
	assign leaf[8890] = f[268] && f[408] && !f[349] && f[606];
	assign leaf[8891] = f[268] && f[408] && f[349] && !f[579];
	assign leaf[8892] = f[268] && f[408] && f[349] && f[579];
	
	// Tree 637, Classifier 7, Iteration: 63
	assign leaf[8893] = !f[372] && !f[405] && !f[492] && !f[205];
	assign leaf[8894] = !f[372] && !f[405] && !f[492] && f[205];
	assign leaf[8895] = !f[372] && !f[405] && f[492] && !f[398];
	assign leaf[8896] = !f[372] && !f[405] && f[492] && f[398];
	assign leaf[8897] = !f[372] && f[405] && !f[346] && !f[435];
	assign leaf[8898] = !f[372] && f[405] && !f[346] && f[435];
	assign leaf[8899] = !f[372] && f[405] && f[346] && !f[316];
	assign leaf[8900] = !f[372] && f[405] && f[346] && f[316];
	assign leaf[8901] = f[372] && !f[460] && !f[318] && !f[349];
	assign leaf[8902] = f[372] && !f[460] && !f[318] && f[349];
	assign leaf[8903] = f[372] && !f[460] && f[318] && !f[516];
	assign leaf[8904] = f[372] && !f[460] && f[318] && f[516];
	assign leaf[8905] = f[372] && f[460] && !f[470] && !f[458];
	assign leaf[8906] = f[372] && f[460] && !f[470] && f[458];
	assign leaf[8907] = f[372] && f[460] && f[470] && !f[577];
	assign leaf[8908] = f[372] && f[460] && f[470] && f[577];
	
	// Tree 638, Classifier 8, Iteration: 63
	assign leaf[8909] = !f[328] && !f[271] && !f[269] && !f[385];
	assign leaf[8910] = !f[328] && !f[271] && !f[269] && f[385];
	assign leaf[8911] = !f[328] && !f[271] && f[269] && !f[326];
	assign leaf[8912] = !f[328] && !f[271] && f[269] && f[326];
	assign leaf[8913] = !f[328] && f[271] && !f[241] && !f[188];
	assign leaf[8914] = !f[328] && f[271] && !f[241] && f[188];
	assign leaf[8915] = !f[328] && f[271] && f[241] && !f[539];
	assign leaf[8916] = !f[328] && f[271] && f[241] && f[539];
	assign leaf[8917] = f[328] && !f[298] && !f[385] && !f[295];
	assign leaf[8918] = f[328] && !f[298] && !f[385] && f[295];
	assign leaf[8919] = f[328] && !f[298] && f[385] && !f[292];
	assign leaf[8920] = f[328] && !f[298] && f[385] && f[292];
	assign leaf[8921] = f[328] && f[298] && !f[240] && !f[356];
	assign leaf[8922] = f[328] && f[298] && !f[240] && f[356];
	assign leaf[8923] = f[328] && f[298] && f[240] && !f[650];
	assign leaf[8924] = f[328] && f[298] && f[240] && f[650];
	
	// Tree 639, Classifier 9, Iteration: 63
	assign leaf[8925] = !f[742] && !f[581] && !f[374] && !f[400];
	assign leaf[8926] = !f[742] && !f[581] && !f[374] && f[400];
	assign leaf[8927] = !f[742] && !f[581] && f[374] && !f[400];
	assign leaf[8928] = !f[742] && !f[581] && f[374] && f[400];
	assign leaf[8929] = !f[742] && f[581] && !f[496] && !f[580];
	assign leaf[8930] = !f[742] && f[581] && !f[496] && f[580];
	assign leaf[8931] = !f[742] && f[581] && f[496] && !f[411];
	assign leaf[8932] = !f[742] && f[581] && f[496] && f[411];
	assign leaf[8933] = f[742] && !f[326] && !f[319] && !f[406];
	assign leaf[8934] = f[742] && !f[326] && !f[319] && f[406];
	assign leaf[8935] = f[742] && !f[326] && f[319];
	assign leaf[8936] = f[742] && f[326] && !f[351] && !f[487];
	assign leaf[8937] = f[742] && f[326] && !f[351] && f[487];
	assign leaf[8938] = f[742] && f[326] && f[351] && !f[660];
	assign leaf[8939] = f[742] && f[326] && f[351] && f[660];
	
	// Tree 640, Classifier 0, Iteration: 64
	assign leaf[8940] = !f[412] && !f[238] && !f[269] && !f[437];
	assign leaf[8941] = !f[412] && !f[238] && !f[269] && f[437];
	assign leaf[8942] = !f[412] && !f[238] && f[269] && !f[354];
	assign leaf[8943] = !f[412] && !f[238] && f[269] && f[354];
	assign leaf[8944] = !f[412] && f[238] && !f[331] && !f[216];
	assign leaf[8945] = !f[412] && f[238] && !f[331] && f[216];
	assign leaf[8946] = !f[412] && f[238] && f[331] && !f[329];
	assign leaf[8947] = !f[412] && f[238] && f[331] && f[329];
	assign leaf[8948] = f[412] && !f[572] && !f[682] && !f[210];
	assign leaf[8949] = f[412] && !f[572] && !f[682] && f[210];
	assign leaf[8950] = f[412] && !f[572] && f[682] && !f[652];
	assign leaf[8951] = f[412] && !f[572] && f[682] && f[652];
	assign leaf[8952] = f[412] && f[572] && !f[321] && !f[387];
	assign leaf[8953] = f[412] && f[572] && !f[321] && f[387];
	assign leaf[8954] = f[412] && f[572] && f[321] && !f[403];
	assign leaf[8955] = f[412] && f[572] && f[321] && f[403];
	
	// Tree 641, Classifier 1, Iteration: 64
	assign leaf[8956] = !f[316] && !f[604] && !f[547] && !f[347];
	assign leaf[8957] = !f[316] && !f[604] && !f[547] && f[347];
	assign leaf[8958] = !f[316] && !f[604] && f[547] && !f[545];
	assign leaf[8959] = !f[316] && !f[604] && f[547] && f[545];
	assign leaf[8960] = !f[316] && f[604] && !f[546] && !f[460];
	assign leaf[8961] = !f[316] && f[604] && !f[546] && f[460];
	assign leaf[8962] = !f[316] && f[604] && f[546] && !f[102];
	assign leaf[8963] = !f[316] && f[604] && f[546] && f[102];
	assign leaf[8964] = f[316] && !f[126];
	assign leaf[8965] = f[316] && f[126];
	
	// Tree 642, Classifier 2, Iteration: 64
	assign leaf[8966] = !f[515] && !f[378] && !f[373] && !f[342];
	assign leaf[8967] = !f[515] && !f[378] && !f[373] && f[342];
	assign leaf[8968] = !f[515] && !f[378] && f[373] && !f[154];
	assign leaf[8969] = !f[515] && !f[378] && f[373] && f[154];
	assign leaf[8970] = !f[515] && f[378] && !f[175] && !f[212];
	assign leaf[8971] = !f[515] && f[378] && !f[175] && f[212];
	assign leaf[8972] = !f[515] && f[378] && f[175] && !f[259];
	assign leaf[8973] = !f[515] && f[378] && f[175] && f[259];
	assign leaf[8974] = f[515] && !f[466] && !f[578] && !f[661];
	assign leaf[8975] = f[515] && !f[466] && !f[578] && f[661];
	assign leaf[8976] = f[515] && !f[466] && f[578] && !f[597];
	assign leaf[8977] = f[515] && !f[466] && f[578] && f[597];
	assign leaf[8978] = f[515] && f[466] && !f[632] && !f[290];
	assign leaf[8979] = f[515] && f[466] && !f[632] && f[290];
	assign leaf[8980] = f[515] && f[466] && f[632] && !f[329];
	assign leaf[8981] = f[515] && f[466] && f[632] && f[329];
	
	// Tree 643, Classifier 3, Iteration: 64
	assign leaf[8982] = !f[346] && !f[290] && !f[292] && !f[376];
	assign leaf[8983] = !f[346] && !f[290] && !f[292] && f[376];
	assign leaf[8984] = !f[346] && !f[290] && f[292] && !f[266];
	assign leaf[8985] = !f[346] && !f[290] && f[292] && f[266];
	assign leaf[8986] = !f[346] && f[290] && !f[320] && !f[129];
	assign leaf[8987] = !f[346] && f[290] && !f[320] && f[129];
	assign leaf[8988] = !f[346] && f[290] && f[320] && !f[238];
	assign leaf[8989] = !f[346] && f[290] && f[320] && f[238];
	assign leaf[8990] = f[346] && !f[321] && !f[403] && !f[327];
	assign leaf[8991] = f[346] && !f[321] && !f[403] && f[327];
	assign leaf[8992] = f[346] && !f[321] && f[403] && !f[636];
	assign leaf[8993] = f[346] && !f[321] && f[403] && f[636];
	assign leaf[8994] = f[346] && f[321] && !f[289] && !f[152];
	assign leaf[8995] = f[346] && f[321] && !f[289] && f[152];
	assign leaf[8996] = f[346] && f[321] && f[289] && !f[627];
	assign leaf[8997] = f[346] && f[321] && f[289] && f[627];
	
	// Tree 644, Classifier 4, Iteration: 64
	assign leaf[8998] = !f[128] && !f[555] && !f[348] && !f[219];
	assign leaf[8999] = !f[128] && !f[555] && !f[348] && f[219];
	assign leaf[9000] = !f[128] && !f[555] && f[348] && !f[716];
	assign leaf[9001] = !f[128] && !f[555] && f[348] && f[716];
	assign leaf[9002] = !f[128] && f[555] && !f[512] && !f[179];
	assign leaf[9003] = !f[128] && f[555] && !f[512] && f[179];
	assign leaf[9004] = !f[128] && f[555] && f[512];
	assign leaf[9005] = f[128] && !f[405] && !f[626] && !f[126];
	assign leaf[9006] = f[128] && !f[405] && !f[626] && f[126];
	assign leaf[9007] = f[128] && !f[405] && f[626];
	assign leaf[9008] = f[128] && f[405] && !f[129];
	assign leaf[9009] = f[128] && f[405] && f[129];
	
	// Tree 645, Classifier 5, Iteration: 64
	assign leaf[9010] = !f[612] && !f[598] && !f[684] && !f[512];
	assign leaf[9011] = !f[612] && !f[598] && !f[684] && f[512];
	assign leaf[9012] = !f[612] && !f[598] && f[684] && !f[576];
	assign leaf[9013] = !f[612] && !f[598] && f[684] && f[576];
	assign leaf[9014] = !f[612] && f[598] && !f[486] && !f[428];
	assign leaf[9015] = !f[612] && f[598] && !f[486] && f[428];
	assign leaf[9016] = !f[612] && f[598] && f[486] && !f[371];
	assign leaf[9017] = !f[612] && f[598] && f[486] && f[371];
	assign leaf[9018] = f[612];
	
	// Tree 646, Classifier 6, Iteration: 64
	assign leaf[9019] = !f[101] && !f[275] && !f[205] && !f[467];
	assign leaf[9020] = !f[101] && !f[275] && !f[205] && f[467];
	assign leaf[9021] = !f[101] && !f[275] && f[205] && !f[182];
	assign leaf[9022] = !f[101] && !f[275] && f[205] && f[182];
	assign leaf[9023] = !f[101] && f[275] && !f[605];
	assign leaf[9024] = !f[101] && f[275] && f[605];
	assign leaf[9025] = f[101] && !f[127] && !f[570];
	assign leaf[9026] = f[101] && !f[127] && f[570] && !f[238];
	assign leaf[9027] = f[101] && !f[127] && f[570] && f[238];
	assign leaf[9028] = f[101] && f[127] && !f[547] && !f[605];
	assign leaf[9029] = f[101] && f[127] && !f[547] && f[605];
	assign leaf[9030] = f[101] && f[127] && f[547] && !f[539];
	assign leaf[9031] = f[101] && f[127] && f[547] && f[539];
	
	// Tree 647, Classifier 7, Iteration: 64
	assign leaf[9032] = !f[325] && !f[205] && !f[542] && !f[314];
	assign leaf[9033] = !f[325] && !f[205] && !f[542] && f[314];
	assign leaf[9034] = !f[325] && !f[205] && f[542] && !f[677];
	assign leaf[9035] = !f[325] && !f[205] && f[542] && f[677];
	assign leaf[9036] = !f[325] && f[205] && !f[605] && !f[575];
	assign leaf[9037] = !f[325] && f[205] && !f[605] && f[575];
	assign leaf[9038] = !f[325] && f[205] && f[605] && !f[263];
	assign leaf[9039] = !f[325] && f[205] && f[605] && f[263];
	assign leaf[9040] = f[325] && !f[150] && !f[437] && !f[548];
	assign leaf[9041] = f[325] && !f[150] && !f[437] && f[548];
	assign leaf[9042] = f[325] && !f[150] && f[437] && !f[176];
	assign leaf[9043] = f[325] && !f[150] && f[437] && f[176];
	assign leaf[9044] = f[325] && f[150] && !f[233] && !f[463];
	assign leaf[9045] = f[325] && f[150] && !f[233] && f[463];
	assign leaf[9046] = f[325] && f[150] && f[233] && !f[430];
	assign leaf[9047] = f[325] && f[150] && f[233] && f[430];
	
	// Tree 648, Classifier 8, Iteration: 64
	assign leaf[9048] = !f[679] && !f[136] && !f[708] && !f[452];
	assign leaf[9049] = !f[679] && !f[136] && !f[708] && f[452];
	assign leaf[9050] = !f[679] && !f[136] && f[708];
	assign leaf[9051] = !f[679] && f[136];
	assign leaf[9052] = f[679] && !f[540] && !f[710] && !f[247];
	assign leaf[9053] = f[679] && !f[540] && !f[710] && f[247];
	assign leaf[9054] = f[679] && !f[540] && f[710];
	assign leaf[9055] = f[679] && f[540] && !f[373] && !f[548];
	assign leaf[9056] = f[679] && f[540] && !f[373] && f[548];
	assign leaf[9057] = f[679] && f[540] && f[373];
	
	// Tree 649, Classifier 9, Iteration: 64
	assign leaf[9058] = !f[717] && !f[718] && !f[128] && !f[517];
	assign leaf[9059] = !f[717] && !f[718] && !f[128] && f[517];
	assign leaf[9060] = !f[717] && !f[718] && f[128] && !f[575];
	assign leaf[9061] = !f[717] && !f[718] && f[128] && f[575];
	assign leaf[9062] = !f[717] && f[718] && !f[488] && !f[318];
	assign leaf[9063] = !f[717] && f[718] && !f[488] && f[318];
	assign leaf[9064] = !f[717] && f[718] && f[488] && !f[287];
	assign leaf[9065] = !f[717] && f[718] && f[488] && f[287];
	assign leaf[9066] = f[717] && !f[211] && !f[299] && !f[238];
	assign leaf[9067] = f[717] && !f[211] && !f[299] && f[238];
	assign leaf[9068] = f[717] && !f[211] && f[299] && !f[231];
	assign leaf[9069] = f[717] && !f[211] && f[299] && f[231];
	assign leaf[9070] = f[717] && f[211] && !f[691] && !f[212];
	assign leaf[9071] = f[717] && f[211] && !f[691] && f[212];
	assign leaf[9072] = f[717] && f[211] && f[691] && !f[438];
	assign leaf[9073] = f[717] && f[211] && f[691] && f[438];
	
	// Tree 650, Classifier 0, Iteration: 65
	assign leaf[9074] = !f[602] && !f[456] && !f[461] && !f[427];
	assign leaf[9075] = !f[602] && !f[456] && !f[461] && f[427];
	assign leaf[9076] = !f[602] && !f[456] && f[461];
	assign leaf[9077] = !f[602] && f[456] && !f[462] && !f[409];
	assign leaf[9078] = !f[602] && f[456] && !f[462] && f[409];
	assign leaf[9079] = !f[602] && f[456] && f[462] && !f[460];
	assign leaf[9080] = !f[602] && f[456] && f[462] && f[460];
	assign leaf[9081] = f[602] && !f[236] && !f[350] && !f[549];
	assign leaf[9082] = f[602] && !f[236] && !f[350] && f[549];
	assign leaf[9083] = f[602] && !f[236] && f[350] && !f[189];
	assign leaf[9084] = f[602] && !f[236] && f[350] && f[189];
	assign leaf[9085] = f[602] && f[236] && !f[463] && !f[483];
	assign leaf[9086] = f[602] && f[236] && !f[463] && f[483];
	assign leaf[9087] = f[602] && f[236] && f[463] && !f[321];
	assign leaf[9088] = f[602] && f[236] && f[463] && f[321];
	
	// Tree 651, Classifier 1, Iteration: 65
	assign leaf[9089] = !f[102] && !f[344] && !f[132] && !f[234];
	assign leaf[9090] = !f[102] && !f[344] && !f[132] && f[234];
	assign leaf[9091] = !f[102] && !f[344] && f[132] && !f[520];
	assign leaf[9092] = !f[102] && !f[344] && f[132] && f[520];
	assign leaf[9093] = !f[102] && f[344] && !f[461];
	assign leaf[9094] = !f[102] && f[344] && f[461];
	assign leaf[9095] = f[102] && !f[629] && !f[626];
	assign leaf[9096] = f[102] && !f[629] && f[626];
	assign leaf[9097] = f[102] && f[629];
	
	// Tree 652, Classifier 2, Iteration: 65
	assign leaf[9098] = !f[154] && !f[133] && !f[219] && !f[213];
	assign leaf[9099] = !f[154] && !f[133] && !f[219] && f[213];
	assign leaf[9100] = !f[154] && !f[133] && f[219] && !f[603];
	assign leaf[9101] = !f[154] && !f[133] && f[219] && f[603];
	assign leaf[9102] = !f[154] && f[133] && !f[156];
	assign leaf[9103] = !f[154] && f[133] && f[156] && !f[351];
	assign leaf[9104] = !f[154] && f[133] && f[156] && f[351];
	assign leaf[9105] = f[154] && !f[625] && !f[290] && !f[486];
	assign leaf[9106] = f[154] && !f[625] && !f[290] && f[486];
	assign leaf[9107] = f[154] && !f[625] && f[290] && !f[299];
	assign leaf[9108] = f[154] && !f[625] && f[290] && f[299];
	assign leaf[9109] = f[154] && f[625] && !f[594] && !f[270];
	assign leaf[9110] = f[154] && f[625] && !f[594] && f[270];
	assign leaf[9111] = f[154] && f[625] && f[594] && !f[346];
	assign leaf[9112] = f[154] && f[625] && f[594] && f[346];
	
	// Tree 653, Classifier 3, Iteration: 65
	assign leaf[9113] = !f[399] && !f[740] && !f[626] && !f[600];
	assign leaf[9114] = !f[399] && !f[740] && !f[626] && f[600];
	assign leaf[9115] = !f[399] && !f[740] && f[626] && !f[629];
	assign leaf[9116] = !f[399] && !f[740] && f[626] && f[629];
	assign leaf[9117] = !f[399] && f[740];
	assign leaf[9118] = f[399] && !f[411] && !f[186] && !f[454];
	assign leaf[9119] = f[399] && !f[411] && !f[186] && f[454];
	assign leaf[9120] = f[399] && !f[411] && f[186] && !f[682];
	assign leaf[9121] = f[399] && !f[411] && f[186] && f[682];
	assign leaf[9122] = f[399] && f[411] && !f[294] && !f[408];
	assign leaf[9123] = f[399] && f[411] && !f[294] && f[408];
	assign leaf[9124] = f[399] && f[411] && f[294] && !f[317];
	assign leaf[9125] = f[399] && f[411] && f[294] && f[317];
	
	// Tree 654, Classifier 4, Iteration: 65
	assign leaf[9126] = !f[744] && !f[121] && !f[102] && !f[656];
	assign leaf[9127] = !f[744] && !f[121] && !f[102] && f[656];
	assign leaf[9128] = !f[744] && !f[121] && f[102] && !f[467];
	assign leaf[9129] = !f[744] && !f[121] && f[102] && f[467];
	assign leaf[9130] = !f[744] && f[121] && !f[484];
	assign leaf[9131] = !f[744] && f[121] && f[484];
	assign leaf[9132] = f[744] && !f[299];
	assign leaf[9133] = f[744] && f[299];
	
	// Tree 655, Classifier 5, Iteration: 65
	assign leaf[9134] = !f[381] && !f[326] && !f[441] && !f[324];
	assign leaf[9135] = !f[381] && !f[326] && !f[441] && f[324];
	assign leaf[9136] = !f[381] && !f[326] && f[441] && !f[661];
	assign leaf[9137] = !f[381] && !f[326] && f[441] && f[661];
	assign leaf[9138] = !f[381] && f[326] && !f[243] && !f[485];
	assign leaf[9139] = !f[381] && f[326] && !f[243] && f[485];
	assign leaf[9140] = !f[381] && f[326] && f[243] && !f[156];
	assign leaf[9141] = !f[381] && f[326] && f[243] && f[156];
	assign leaf[9142] = f[381] && !f[327] && !f[132] && !f[244];
	assign leaf[9143] = f[381] && !f[327] && !f[132] && f[244];
	assign leaf[9144] = f[381] && !f[327] && f[132] && !f[243];
	assign leaf[9145] = f[381] && !f[327] && f[132] && f[243];
	assign leaf[9146] = f[381] && f[327] && !f[294] && !f[409];
	assign leaf[9147] = f[381] && f[327] && !f[294] && f[409];
	assign leaf[9148] = f[381] && f[327] && f[294] && !f[653];
	assign leaf[9149] = f[381] && f[327] && f[294] && f[653];
	
	// Tree 656, Classifier 6, Iteration: 65
	assign leaf[9150] = !f[268] && !f[136] && !f[231] && !f[636];
	assign leaf[9151] = !f[268] && !f[136] && !f[231] && f[636];
	assign leaf[9152] = !f[268] && !f[136] && f[231] && !f[347];
	assign leaf[9153] = !f[268] && !f[136] && f[231] && f[347];
	assign leaf[9154] = !f[268] && f[136];
	assign leaf[9155] = f[268] && !f[380] && !f[570] && !f[512];
	assign leaf[9156] = f[268] && !f[380] && !f[570] && f[512];
	assign leaf[9157] = f[268] && !f[380] && f[570] && !f[490];
	assign leaf[9158] = f[268] && !f[380] && f[570] && f[490];
	assign leaf[9159] = f[268] && f[380] && !f[324] && !f[486];
	assign leaf[9160] = f[268] && f[380] && !f[324] && f[486];
	assign leaf[9161] = f[268] && f[380] && f[324] && !f[161];
	assign leaf[9162] = f[268] && f[380] && f[324] && f[161];
	
	// Tree 657, Classifier 7, Iteration: 65
	assign leaf[9163] = !f[269] && !f[601] && !f[684] && !f[545];
	assign leaf[9164] = !f[269] && !f[601] && !f[684] && f[545];
	assign leaf[9165] = !f[269] && !f[601] && f[684] && !f[660];
	assign leaf[9166] = !f[269] && !f[601] && f[684] && f[660];
	assign leaf[9167] = !f[269] && f[601] && !f[177] && !f[453];
	assign leaf[9168] = !f[269] && f[601] && !f[177] && f[453];
	assign leaf[9169] = !f[269] && f[601] && f[177] && !f[550];
	assign leaf[9170] = !f[269] && f[601] && f[177] && f[550];
	assign leaf[9171] = f[269] && !f[577] && !f[663] && !f[482];
	assign leaf[9172] = f[269] && !f[577] && !f[663] && f[482];
	assign leaf[9173] = f[269] && !f[577] && f[663] && !f[291];
	assign leaf[9174] = f[269] && !f[577] && f[663] && f[291];
	assign leaf[9175] = f[269] && f[577] && !f[522] && !f[465];
	assign leaf[9176] = f[269] && f[577] && !f[522] && f[465];
	assign leaf[9177] = f[269] && f[577] && f[522] && !f[660];
	assign leaf[9178] = f[269] && f[577] && f[522] && f[660];
	
	// Tree 658, Classifier 8, Iteration: 65
	assign leaf[9179] = !f[341] && !f[491] && !f[294] && !f[303];
	assign leaf[9180] = !f[341] && !f[491] && !f[294] && f[303];
	assign leaf[9181] = !f[341] && !f[491] && f[294] && !f[380];
	assign leaf[9182] = !f[341] && !f[491] && f[294] && f[380];
	assign leaf[9183] = !f[341] && f[491] && !f[436] && !f[494];
	assign leaf[9184] = !f[341] && f[491] && !f[436] && f[494];
	assign leaf[9185] = !f[341] && f[491] && f[436] && !f[352];
	assign leaf[9186] = !f[341] && f[491] && f[436] && f[352];
	assign leaf[9187] = f[341] && !f[315] && !f[662];
	assign leaf[9188] = f[341] && !f[315] && f[662];
	assign leaf[9189] = f[341] && f[315] && !f[464] && !f[486];
	assign leaf[9190] = f[341] && f[315] && !f[464] && f[486];
	assign leaf[9191] = f[341] && f[315] && f[464] && !f[601];
	assign leaf[9192] = f[341] && f[315] && f[464] && f[601];
	
	// Tree 659, Classifier 9, Iteration: 65
	assign leaf[9193] = !f[687] && !f[509] && !f[584] && !f[320];
	assign leaf[9194] = !f[687] && !f[509] && !f[584] && f[320];
	assign leaf[9195] = !f[687] && !f[509] && f[584];
	assign leaf[9196] = !f[687] && f[509] && !f[236];
	assign leaf[9197] = !f[687] && f[509] && f[236] && !f[662];
	assign leaf[9198] = !f[687] && f[509] && f[236] && f[662];
	assign leaf[9199] = f[687] && !f[573] && !f[378] && !f[489];
	assign leaf[9200] = f[687] && !f[573] && !f[378] && f[489];
	assign leaf[9201] = f[687] && !f[573] && f[378] && !f[352];
	assign leaf[9202] = f[687] && !f[573] && f[378] && f[352];
	assign leaf[9203] = f[687] && f[573] && !f[158] && !f[484];
	assign leaf[9204] = f[687] && f[573] && !f[158] && f[484];
	assign leaf[9205] = f[687] && f[573] && f[158] && !f[428];
	assign leaf[9206] = f[687] && f[573] && f[158] && f[428];
	
	// Tree 660, Classifier 0, Iteration: 66
	assign leaf[9207] = !f[572] && !f[684] && !f[541] && !f[629];
	assign leaf[9208] = !f[572] && !f[684] && !f[541] && f[629];
	assign leaf[9209] = !f[572] && !f[684] && f[541] && !f[212];
	assign leaf[9210] = !f[572] && !f[684] && f[541] && f[212];
	assign leaf[9211] = !f[572] && f[684] && !f[574] && !f[353];
	assign leaf[9212] = !f[572] && f[684] && !f[574] && f[353];
	assign leaf[9213] = !f[572] && f[684] && f[574] && !f[596];
	assign leaf[9214] = !f[572] && f[684] && f[574] && f[596];
	assign leaf[9215] = f[572] && !f[683] && !f[598] && !f[319];
	assign leaf[9216] = f[572] && !f[683] && !f[598] && f[319];
	assign leaf[9217] = f[572] && !f[683] && f[598] && !f[608];
	assign leaf[9218] = f[572] && !f[683] && f[598] && f[608];
	assign leaf[9219] = f[572] && f[683] && !f[548];
	assign leaf[9220] = f[572] && f[683] && f[548];
	
	// Tree 661, Classifier 1, Iteration: 66
	assign leaf[9221] = !f[556] && !f[511] && !f[323] && !f[183];
	assign leaf[9222] = !f[556] && !f[511] && !f[323] && f[183];
	assign leaf[9223] = !f[556] && !f[511] && f[323] && !f[351];
	assign leaf[9224] = !f[556] && !f[511] && f[323] && f[351];
	assign leaf[9225] = !f[556] && f[511] && !f[622];
	assign leaf[9226] = !f[556] && f[511] && f[622];
	assign leaf[9227] = f[556];
	
	// Tree 662, Classifier 2, Iteration: 66
	assign leaf[9228] = !f[242] && !f[183] && !f[326] && !f[240];
	assign leaf[9229] = !f[242] && !f[183] && !f[326] && f[240];
	assign leaf[9230] = !f[242] && !f[183] && f[326] && !f[269];
	assign leaf[9231] = !f[242] && !f[183] && f[326] && f[269];
	assign leaf[9232] = !f[242] && f[183] && !f[240] && !f[188];
	assign leaf[9233] = !f[242] && f[183] && !f[240] && f[188];
	assign leaf[9234] = !f[242] && f[183] && f[240] && !f[500];
	assign leaf[9235] = !f[242] && f[183] && f[240] && f[500];
	assign leaf[9236] = f[242] && !f[184] && !f[129] && !f[324];
	assign leaf[9237] = f[242] && !f[184] && !f[129] && f[324];
	assign leaf[9238] = f[242] && !f[184] && f[129] && !f[238];
	assign leaf[9239] = f[242] && !f[184] && f[129] && f[238];
	assign leaf[9240] = f[242] && f[184] && !f[540] && !f[688];
	assign leaf[9241] = f[242] && f[184] && !f[540] && f[688];
	assign leaf[9242] = f[242] && f[184] && f[540] && !f[651];
	assign leaf[9243] = f[242] && f[184] && f[540] && f[651];
	
	// Tree 663, Classifier 3, Iteration: 66
	assign leaf[9244] = !f[429] && !f[213] && !f[713] && !f[458];
	assign leaf[9245] = !f[429] && !f[213] && !f[713] && f[458];
	assign leaf[9246] = !f[429] && !f[213] && f[713] && !f[323];
	assign leaf[9247] = !f[429] && !f[213] && f[713] && f[323];
	assign leaf[9248] = !f[429] && f[213] && !f[126] && !f[570];
	assign leaf[9249] = !f[429] && f[213] && !f[126] && f[570];
	assign leaf[9250] = !f[429] && f[213] && f[126] && !f[487];
	assign leaf[9251] = !f[429] && f[213] && f[126] && f[487];
	assign leaf[9252] = f[429] && !f[459] && !f[483] && !f[485];
	assign leaf[9253] = f[429] && !f[459] && !f[483] && f[485];
	assign leaf[9254] = f[429] && !f[459] && f[483] && !f[498];
	assign leaf[9255] = f[429] && !f[459] && f[483] && f[498];
	assign leaf[9256] = f[429] && f[459] && !f[346] && !f[580];
	assign leaf[9257] = f[429] && f[459] && !f[346] && f[580];
	assign leaf[9258] = f[429] && f[459] && f[346] && !f[182];
	assign leaf[9259] = f[429] && f[459] && f[346] && f[182];
	
	// Tree 664, Classifier 4, Iteration: 66
	assign leaf[9260] = !f[738] && !f[96] && !f[747] && !f[384];
	assign leaf[9261] = !f[738] && !f[96] && !f[747] && f[384];
	assign leaf[9262] = !f[738] && !f[96] && f[747];
	assign leaf[9263] = !f[738] && f[96];
	assign leaf[9264] = f[738] && !f[269];
	assign leaf[9265] = f[738] && f[269];
	
	// Tree 665, Classifier 5, Iteration: 66
	assign leaf[9266] = !f[99] && !f[188] && !f[244] && !f[239];
	assign leaf[9267] = !f[99] && !f[188] && !f[244] && f[239];
	assign leaf[9268] = !f[99] && !f[188] && f[244] && !f[267];
	assign leaf[9269] = !f[99] && !f[188] && f[244] && f[267];
	assign leaf[9270] = !f[99] && f[188] && !f[273] && !f[271];
	assign leaf[9271] = !f[99] && f[188] && !f[273] && f[271];
	assign leaf[9272] = !f[99] && f[188] && f[273] && !f[269];
	assign leaf[9273] = !f[99] && f[188] && f[273] && f[269];
	assign leaf[9274] = f[99] && !f[240] && !f[431] && !f[344];
	assign leaf[9275] = f[99] && !f[240] && !f[431] && f[344];
	assign leaf[9276] = f[99] && !f[240] && f[431] && !f[317];
	assign leaf[9277] = f[99] && !f[240] && f[431] && f[317];
	assign leaf[9278] = f[99] && f[240] && !f[185];
	assign leaf[9279] = f[99] && f[240] && f[185];
	
	// Tree 666, Classifier 6, Iteration: 66
	assign leaf[9280] = !f[91] && !f[213] && !f[324] && !f[323];
	assign leaf[9281] = !f[91] && !f[213] && !f[324] && f[323];
	assign leaf[9282] = !f[91] && !f[213] && f[324] && !f[238];
	assign leaf[9283] = !f[91] && !f[213] && f[324] && f[238];
	assign leaf[9284] = !f[91] && f[213] && !f[325] && !f[356];
	assign leaf[9285] = !f[91] && f[213] && !f[325] && f[356];
	assign leaf[9286] = !f[91] && f[213] && f[325] && !f[190];
	assign leaf[9287] = !f[91] && f[213] && f[325] && f[190];
	assign leaf[9288] = f[91];
	
	// Tree 667, Classifier 7, Iteration: 66
	assign leaf[9289] = !f[129] && !f[148] && !f[160] && !f[150];
	assign leaf[9290] = !f[129] && !f[148] && !f[160] && f[150];
	assign leaf[9291] = !f[129] && !f[148] && f[160];
	assign leaf[9292] = !f[129] && f[148] && !f[153] && !f[146];
	assign leaf[9293] = !f[129] && f[148] && !f[153] && f[146];
	assign leaf[9294] = !f[129] && f[148] && f[153] && !f[520];
	assign leaf[9295] = !f[129] && f[148] && f[153] && f[520];
	assign leaf[9296] = f[129];
	
	// Tree 668, Classifier 8, Iteration: 66
	assign leaf[9297] = !f[465] && !f[520] && !f[207] && !f[627];
	assign leaf[9298] = !f[465] && !f[520] && !f[207] && f[627];
	assign leaf[9299] = !f[465] && !f[520] && f[207] && !f[600];
	assign leaf[9300] = !f[465] && !f[520] && f[207] && f[600];
	assign leaf[9301] = !f[465] && f[520] && !f[434] && !f[602];
	assign leaf[9302] = !f[465] && f[520] && !f[434] && f[602];
	assign leaf[9303] = !f[465] && f[520] && f[434] && !f[235];
	assign leaf[9304] = !f[465] && f[520] && f[434] && f[235];
	assign leaf[9305] = f[465] && !f[151] && !f[216] && !f[266];
	assign leaf[9306] = f[465] && !f[151] && !f[216] && f[266];
	assign leaf[9307] = f[465] && !f[151] && f[216] && !f[125];
	assign leaf[9308] = f[465] && !f[151] && f[216] && f[125];
	assign leaf[9309] = f[465] && f[151] && !f[487] && !f[313];
	assign leaf[9310] = f[465] && f[151] && !f[487] && f[313];
	assign leaf[9311] = f[465] && f[151] && f[487] && !f[543];
	assign leaf[9312] = f[465] && f[151] && f[487] && f[543];
	
	// Tree 669, Classifier 9, Iteration: 66
	assign leaf[9313] = !f[368] && !f[498] && !f[184] && !f[240];
	assign leaf[9314] = !f[368] && !f[498] && !f[184] && f[240];
	assign leaf[9315] = !f[368] && !f[498] && f[184] && !f[240];
	assign leaf[9316] = !f[368] && !f[498] && f[184] && f[240];
	assign leaf[9317] = !f[368] && f[498] && !f[584] && !f[682];
	assign leaf[9318] = !f[368] && f[498] && !f[584] && f[682];
	assign leaf[9319] = !f[368] && f[498] && f[584];
	assign leaf[9320] = f[368] && !f[347] && !f[385] && !f[520];
	assign leaf[9321] = f[368] && !f[347] && !f[385] && f[520];
	assign leaf[9322] = f[368] && !f[347] && f[385] && !f[398];
	assign leaf[9323] = f[368] && !f[347] && f[385] && f[398];
	assign leaf[9324] = f[368] && f[347] && !f[320];
	assign leaf[9325] = f[368] && f[347] && f[320];
	
	// Tree 670, Classifier 0, Iteration: 67
	assign leaf[9326] = !f[444] && !f[633] && !f[580] && !f[713];
	assign leaf[9327] = !f[444] && !f[633] && !f[580] && f[713];
	assign leaf[9328] = !f[444] && !f[633] && f[580] && !f[354];
	assign leaf[9329] = !f[444] && !f[633] && f[580] && f[354];
	assign leaf[9330] = !f[444] && f[633] && !f[552] && !f[658];
	assign leaf[9331] = !f[444] && f[633] && !f[552] && f[658];
	assign leaf[9332] = !f[444] && f[633] && f[552] && !f[544];
	assign leaf[9333] = !f[444] && f[633] && f[552] && f[544];
	assign leaf[9334] = f[444] && !f[152] && !f[317];
	assign leaf[9335] = f[444] && !f[152] && f[317];
	assign leaf[9336] = f[444] && f[152];
	
	// Tree 671, Classifier 1, Iteration: 67
	assign leaf[9337] = !f[378] && !f[322] && !f[517] && !f[434];
	assign leaf[9338] = !f[378] && !f[322] && !f[517] && f[434];
	assign leaf[9339] = !f[378] && !f[322] && f[517] && !f[549];
	assign leaf[9340] = !f[378] && !f[322] && f[517] && f[549];
	assign leaf[9341] = !f[378] && f[322] && !f[434] && !f[292];
	assign leaf[9342] = !f[378] && f[322] && !f[434] && f[292];
	assign leaf[9343] = !f[378] && f[322] && f[434] && !f[292];
	assign leaf[9344] = !f[378] && f[322] && f[434] && f[292];
	assign leaf[9345] = f[378] && !f[294] && !f[182] && !f[574];
	assign leaf[9346] = f[378] && !f[294] && !f[182] && f[574];
	assign leaf[9347] = f[378] && !f[294] && f[182] && !f[579];
	assign leaf[9348] = f[378] && !f[294] && f[182] && f[579];
	assign leaf[9349] = f[378] && f[294] && !f[375] && !f[596];
	assign leaf[9350] = f[378] && f[294] && !f[375] && f[596];
	assign leaf[9351] = f[378] && f[294] && f[375] && !f[657];
	assign leaf[9352] = f[378] && f[294] && f[375] && f[657];
	
	// Tree 672, Classifier 2, Iteration: 67
	assign leaf[9353] = !f[485] && !f[403] && !f[512] && !f[257];
	assign leaf[9354] = !f[485] && !f[403] && !f[512] && f[257];
	assign leaf[9355] = !f[485] && !f[403] && f[512] && !f[459];
	assign leaf[9356] = !f[485] && !f[403] && f[512] && f[459];
	assign leaf[9357] = !f[485] && f[403] && !f[428] && !f[122];
	assign leaf[9358] = !f[485] && f[403] && !f[428] && f[122];
	assign leaf[9359] = !f[485] && f[403] && f[428] && !f[294];
	assign leaf[9360] = !f[485] && f[403] && f[428] && f[294];
	assign leaf[9361] = f[485] && !f[690] && !f[685] && !f[433];
	assign leaf[9362] = f[485] && !f[690] && !f[685] && f[433];
	assign leaf[9363] = f[485] && !f[690] && f[685] && !f[607];
	assign leaf[9364] = f[485] && !f[690] && f[685] && f[607];
	assign leaf[9365] = f[485] && f[690] && !f[187];
	assign leaf[9366] = f[485] && f[690] && f[187];
	
	// Tree 673, Classifier 3, Iteration: 67
	assign leaf[9367] = !f[386] && !f[537] && !f[570] && !f[460];
	assign leaf[9368] = !f[386] && !f[537] && !f[570] && f[460];
	assign leaf[9369] = !f[386] && !f[537] && f[570] && !f[600];
	assign leaf[9370] = !f[386] && !f[537] && f[570] && f[600];
	assign leaf[9371] = !f[386] && f[537] && !f[302] && !f[602];
	assign leaf[9372] = !f[386] && f[537] && !f[302] && f[602];
	assign leaf[9373] = !f[386] && f[537] && f[302] && !f[483];
	assign leaf[9374] = !f[386] && f[537] && f[302] && f[483];
	assign leaf[9375] = f[386] && !f[355];
	assign leaf[9376] = f[386] && f[355] && !f[580] && !f[185];
	assign leaf[9377] = f[386] && f[355] && !f[580] && f[185];
	assign leaf[9378] = f[386] && f[355] && f[580] && !f[259];
	assign leaf[9379] = f[386] && f[355] && f[580] && f[259];
	
	// Tree 674, Classifier 4, Iteration: 67
	assign leaf[9380] = !f[429] && !f[349] && !f[237] && !f[293];
	assign leaf[9381] = !f[429] && !f[349] && !f[237] && f[293];
	assign leaf[9382] = !f[429] && !f[349] && f[237] && !f[211];
	assign leaf[9383] = !f[429] && !f[349] && f[237] && f[211];
	assign leaf[9384] = !f[429] && f[349] && !f[467] && !f[454];
	assign leaf[9385] = !f[429] && f[349] && !f[467] && f[454];
	assign leaf[9386] = !f[429] && f[349] && f[467] && !f[184];
	assign leaf[9387] = !f[429] && f[349] && f[467] && f[184];
	assign leaf[9388] = f[429] && !f[205] && !f[214] && !f[210];
	assign leaf[9389] = f[429] && !f[205] && !f[214] && f[210];
	assign leaf[9390] = f[429] && !f[205] && f[214] && !f[272];
	assign leaf[9391] = f[429] && !f[205] && f[214] && f[272];
	assign leaf[9392] = f[429] && f[205] && !f[289] && !f[413];
	assign leaf[9393] = f[429] && f[205] && !f[289] && f[413];
	assign leaf[9394] = f[429] && f[205] && f[289] && !f[265];
	assign leaf[9395] = f[429] && f[205] && f[289] && f[265];
	
	// Tree 675, Classifier 5, Iteration: 67
	assign leaf[9396] = !f[200] && !f[436] && !f[485] && !f[292];
	assign leaf[9397] = !f[200] && !f[436] && !f[485] && f[292];
	assign leaf[9398] = !f[200] && !f[436] && f[485] && !f[352];
	assign leaf[9399] = !f[200] && !f[436] && f[485] && f[352];
	assign leaf[9400] = !f[200] && f[436] && !f[354] && !f[384];
	assign leaf[9401] = !f[200] && f[436] && !f[354] && f[384];
	assign leaf[9402] = !f[200] && f[436] && f[354] && !f[324];
	assign leaf[9403] = !f[200] && f[436] && f[354] && f[324];
	assign leaf[9404] = f[200];
	
	// Tree 676, Classifier 6, Iteration: 67
	assign leaf[9405] = !f[602] && !f[126] && !f[629] && !f[291];
	assign leaf[9406] = !f[602] && !f[126] && !f[629] && f[291];
	assign leaf[9407] = !f[602] && !f[126] && f[629] && !f[522];
	assign leaf[9408] = !f[602] && !f[126] && f[629] && f[522];
	assign leaf[9409] = !f[602] && f[126] && !f[574] && !f[491];
	assign leaf[9410] = !f[602] && f[126] && !f[574] && f[491];
	assign leaf[9411] = !f[602] && f[126] && f[574] && !f[208];
	assign leaf[9412] = !f[602] && f[126] && f[574] && f[208];
	assign leaf[9413] = f[602] && !f[486] && !f[543] && !f[544];
	assign leaf[9414] = f[602] && !f[486] && !f[543] && f[544];
	assign leaf[9415] = f[602] && !f[486] && f[543] && !f[426];
	assign leaf[9416] = f[602] && !f[486] && f[543] && f[426];
	assign leaf[9417] = f[602] && f[486] && !f[189] && !f[374];
	assign leaf[9418] = f[602] && f[486] && !f[189] && f[374];
	assign leaf[9419] = f[602] && f[486] && f[189] && !f[521];
	assign leaf[9420] = f[602] && f[486] && f[189] && f[521];
	
	// Tree 677, Classifier 7, Iteration: 67
	assign leaf[9421] = !f[473] && !f[441] && !f[206] && !f[432];
	assign leaf[9422] = !f[473] && !f[441] && !f[206] && f[432];
	assign leaf[9423] = !f[473] && !f[441] && f[206] && !f[260];
	assign leaf[9424] = !f[473] && !f[441] && f[206] && f[260];
	assign leaf[9425] = !f[473] && f[441] && !f[542] && !f[241];
	assign leaf[9426] = !f[473] && f[441] && !f[542] && f[241];
	assign leaf[9427] = !f[473] && f[441] && f[542] && !f[651];
	assign leaf[9428] = !f[473] && f[441] && f[542] && f[651];
	assign leaf[9429] = f[473];
	
	// Tree 678, Classifier 8, Iteration: 67
	assign leaf[9430] = !f[382] && !f[326] && !f[263] && !f[290];
	assign leaf[9431] = !f[382] && !f[326] && !f[263] && f[290];
	assign leaf[9432] = !f[382] && !f[326] && f[263] && !f[296];
	assign leaf[9433] = !f[382] && !f[326] && f[263] && f[296];
	assign leaf[9434] = !f[382] && f[326] && !f[215] && !f[356];
	assign leaf[9435] = !f[382] && f[326] && !f[215] && f[356];
	assign leaf[9436] = !f[382] && f[326] && f[215] && !f[296];
	assign leaf[9437] = !f[382] && f[326] && f[215] && f[296];
	assign leaf[9438] = f[382] && !f[352] && !f[494] && !f[685];
	assign leaf[9439] = f[382] && !f[352] && !f[494] && f[685];
	assign leaf[9440] = f[382] && !f[352] && f[494] && !f[411];
	assign leaf[9441] = f[382] && !f[352] && f[494] && f[411];
	assign leaf[9442] = f[382] && f[352] && !f[483] && !f[513];
	assign leaf[9443] = f[382] && f[352] && !f[483] && f[513];
	assign leaf[9444] = f[382] && f[352] && f[483] && !f[625];
	assign leaf[9445] = f[382] && f[352] && f[483] && f[625];
	
	// Tree 679, Classifier 9, Iteration: 67
	assign leaf[9446] = !f[351] && !f[383] && !f[381] && !f[519];
	assign leaf[9447] = !f[351] && !f[383] && !f[381] && f[519];
	assign leaf[9448] = !f[351] && !f[383] && f[381] && !f[270];
	assign leaf[9449] = !f[351] && !f[383] && f[381] && f[270];
	assign leaf[9450] = !f[351] && f[383] && !f[407] && !f[291];
	assign leaf[9451] = !f[351] && f[383] && !f[407] && f[291];
	assign leaf[9452] = !f[351] && f[383] && f[407] && !f[349];
	assign leaf[9453] = !f[351] && f[383] && f[407] && f[349];
	assign leaf[9454] = f[351] && !f[326] && !f[382] && !f[438];
	assign leaf[9455] = f[351] && !f[326] && !f[382] && f[438];
	assign leaf[9456] = f[351] && !f[326] && f[382] && !f[466];
	assign leaf[9457] = f[351] && !f[326] && f[382] && f[466];
	assign leaf[9458] = f[351] && f[326] && !f[213] && !f[600];
	assign leaf[9459] = f[351] && f[326] && !f[213] && f[600];
	assign leaf[9460] = f[351] && f[326] && f[213] && !f[538];
	assign leaf[9461] = f[351] && f[326] && f[213] && f[538];
	
	// Tree 680, Classifier 0, Iteration: 68
	assign leaf[9462] = !f[444] && !f[516] && !f[379] && !f[486];
	assign leaf[9463] = !f[444] && !f[516] && !f[379] && f[486];
	assign leaf[9464] = !f[444] && !f[516] && f[379] && !f[268];
	assign leaf[9465] = !f[444] && !f[516] && f[379] && f[268];
	assign leaf[9466] = !f[444] && f[516] && !f[437] && !f[206];
	assign leaf[9467] = !f[444] && f[516] && !f[437] && f[206];
	assign leaf[9468] = !f[444] && f[516] && f[437] && !f[596];
	assign leaf[9469] = !f[444] && f[516] && f[437] && f[596];
	assign leaf[9470] = f[444] && !f[514] && !f[357];
	assign leaf[9471] = f[444] && !f[514] && f[357];
	assign leaf[9472] = f[444] && f[514] && !f[602];
	assign leaf[9473] = f[444] && f[514] && f[602];
	
	// Tree 681, Classifier 1, Iteration: 68
	assign leaf[9474] = !f[606] && !f[204] && !f[661] && !f[263];
	assign leaf[9475] = !f[606] && !f[204] && !f[661] && f[263];
	assign leaf[9476] = !f[606] && !f[204] && f[661] && !f[208];
	assign leaf[9477] = !f[606] && !f[204] && f[661] && f[208];
	assign leaf[9478] = !f[606] && f[204] && !f[321];
	assign leaf[9479] = !f[606] && f[204] && f[321];
	assign leaf[9480] = f[606] && !f[267] && !f[488] && !f[547];
	assign leaf[9481] = f[606] && !f[267] && !f[488] && f[547];
	assign leaf[9482] = f[606] && !f[267] && f[488];
	assign leaf[9483] = f[606] && f[267] && !f[149] && !f[661];
	assign leaf[9484] = f[606] && f[267] && !f[149] && f[661];
	assign leaf[9485] = f[606] && f[267] && f[149];
	
	// Tree 682, Classifier 2, Iteration: 68
	assign leaf[9486] = !f[323] && !f[261] && !f[292] && !f[399];
	assign leaf[9487] = !f[323] && !f[261] && !f[292] && f[399];
	assign leaf[9488] = !f[323] && !f[261] && f[292] && !f[322];
	assign leaf[9489] = !f[323] && !f[261] && f[292] && f[322];
	assign leaf[9490] = !f[323] && f[261] && !f[285] && !f[625];
	assign leaf[9491] = !f[323] && f[261] && !f[285] && f[625];
	assign leaf[9492] = !f[323] && f[261] && f[285] && !f[484];
	assign leaf[9493] = !f[323] && f[261] && f[285] && f[484];
	assign leaf[9494] = f[323] && !f[217] && !f[528] && !f[439];
	assign leaf[9495] = f[323] && !f[217] && !f[528] && f[439];
	assign leaf[9496] = f[323] && !f[217] && f[528] && !f[567];
	assign leaf[9497] = f[323] && !f[217] && f[528] && f[567];
	assign leaf[9498] = f[323] && f[217] && !f[607] && !f[508];
	assign leaf[9499] = f[323] && f[217] && !f[607] && f[508];
	assign leaf[9500] = f[323] && f[217] && f[607] && !f[511];
	assign leaf[9501] = f[323] && f[217] && f[607] && f[511];
	
	// Tree 683, Classifier 3, Iteration: 68
	assign leaf[9502] = !f[682] && !f[626] && !f[602] && !f[714];
	assign leaf[9503] = !f[682] && !f[626] && !f[602] && f[714];
	assign leaf[9504] = !f[682] && !f[626] && f[602] && !f[598];
	assign leaf[9505] = !f[682] && !f[626] && f[602] && f[598];
	assign leaf[9506] = !f[682] && f[626] && !f[431] && !f[207];
	assign leaf[9507] = !f[682] && f[626] && !f[431] && f[207];
	assign leaf[9508] = !f[682] && f[626] && f[431] && !f[485];
	assign leaf[9509] = !f[682] && f[626] && f[431] && f[485];
	assign leaf[9510] = f[682] && !f[541] && !f[320] && !f[602];
	assign leaf[9511] = f[682] && !f[541] && !f[320] && f[602];
	assign leaf[9512] = f[682] && !f[541] && f[320] && !f[598];
	assign leaf[9513] = f[682] && !f[541] && f[320] && f[598];
	assign leaf[9514] = f[682] && f[541] && !f[514] && !f[299];
	assign leaf[9515] = f[682] && f[541] && !f[514] && f[299];
	assign leaf[9516] = f[682] && f[541] && f[514] && !f[407];
	assign leaf[9517] = f[682] && f[541] && f[514] && f[407];
	
	// Tree 684, Classifier 4, Iteration: 68
	assign leaf[9518] = !f[179] && !f[690] && !f[525] && !f[539];
	assign leaf[9519] = !f[179] && !f[690] && !f[525] && f[539];
	assign leaf[9520] = !f[179] && !f[690] && f[525] && !f[596];
	assign leaf[9521] = !f[179] && !f[690] && f[525] && f[596];
	assign leaf[9522] = !f[179] && f[690] && !f[236] && !f[239];
	assign leaf[9523] = !f[179] && f[690] && !f[236] && f[239];
	assign leaf[9524] = !f[179] && f[690] && f[236] && !f[181];
	assign leaf[9525] = !f[179] && f[690] && f[236] && f[181];
	assign leaf[9526] = f[179] && !f[263] && !f[152] && !f[181];
	assign leaf[9527] = f[179] && !f[263] && !f[152] && f[181];
	assign leaf[9528] = f[179] && !f[263] && f[152] && !f[483];
	assign leaf[9529] = f[179] && !f[263] && f[152] && f[483];
	assign leaf[9530] = f[179] && f[263] && !f[213] && !f[354];
	assign leaf[9531] = f[179] && f[263] && !f[213] && f[354];
	assign leaf[9532] = f[179] && f[263] && f[213] && !f[182];
	assign leaf[9533] = f[179] && f[263] && f[213] && f[182];
	
	// Tree 685, Classifier 5, Iteration: 68
	assign leaf[9534] = !f[120] && !f[686] && !f[598] && !f[509];
	assign leaf[9535] = !f[120] && !f[686] && !f[598] && f[509];
	assign leaf[9536] = !f[120] && !f[686] && f[598] && !f[214];
	assign leaf[9537] = !f[120] && !f[686] && f[598] && f[214];
	assign leaf[9538] = !f[120] && f[686] && !f[546] && !f[345];
	assign leaf[9539] = !f[120] && f[686] && !f[546] && f[345];
	assign leaf[9540] = !f[120] && f[686] && f[546] && !f[682];
	assign leaf[9541] = !f[120] && f[686] && f[546] && f[682];
	assign leaf[9542] = f[120] && !f[204] && !f[553];
	assign leaf[9543] = f[120] && !f[204] && f[553];
	assign leaf[9544] = f[120] && f[204];
	
	// Tree 686, Classifier 6, Iteration: 68
	assign leaf[9545] = !f[270] && !f[514] && !f[406] && !f[267];
	assign leaf[9546] = !f[270] && !f[514] && !f[406] && f[267];
	assign leaf[9547] = !f[270] && !f[514] && f[406] && !f[462];
	assign leaf[9548] = !f[270] && !f[514] && f[406] && f[462];
	assign leaf[9549] = !f[270] && f[514] && !f[401] && !f[153];
	assign leaf[9550] = !f[270] && f[514] && !f[401] && f[153];
	assign leaf[9551] = !f[270] && f[514] && f[401] && !f[571];
	assign leaf[9552] = !f[270] && f[514] && f[401] && f[571];
	assign leaf[9553] = f[270] && !f[272] && !f[541] && !f[325];
	assign leaf[9554] = f[270] && !f[272] && !f[541] && f[325];
	assign leaf[9555] = f[270] && !f[272] && f[541] && !f[540];
	assign leaf[9556] = f[270] && !f[272] && f[541] && f[540];
	assign leaf[9557] = f[270] && f[272] && !f[186] && !f[355];
	assign leaf[9558] = f[270] && f[272] && !f[186] && f[355];
	assign leaf[9559] = f[270] && f[272] && f[186] && !f[468];
	assign leaf[9560] = f[270] && f[272] && f[186] && f[468];
	
	// Tree 687, Classifier 7, Iteration: 68
	assign leaf[9561] = !f[528] && !f[510] && !f[527] && !f[274];
	assign leaf[9562] = !f[528] && !f[510] && !f[527] && f[274];
	assign leaf[9563] = !f[528] && !f[510] && f[527] && !f[242];
	assign leaf[9564] = !f[528] && !f[510] && f[527] && f[242];
	assign leaf[9565] = !f[528] && f[510] && !f[660] && !f[656];
	assign leaf[9566] = !f[528] && f[510] && !f[660] && f[656];
	assign leaf[9567] = !f[528] && f[510] && f[660] && !f[457];
	assign leaf[9568] = !f[528] && f[510] && f[660] && f[457];
	assign leaf[9569] = f[528] && !f[353];
	assign leaf[9570] = f[528] && f[353];
	
	// Tree 688, Classifier 8, Iteration: 68
	assign leaf[9571] = !f[314] && !f[290] && !f[316] && !f[232];
	assign leaf[9572] = !f[314] && !f[290] && !f[316] && f[232];
	assign leaf[9573] = !f[314] && !f[290] && f[316] && !f[234];
	assign leaf[9574] = !f[314] && !f[290] && f[316] && f[234];
	assign leaf[9575] = !f[314] && f[290] && !f[348] && !f[544];
	assign leaf[9576] = !f[314] && f[290] && !f[348] && f[544];
	assign leaf[9577] = !f[314] && f[290] && f[348] && !f[373];
	assign leaf[9578] = !f[314] && f[290] && f[348] && f[373];
	assign leaf[9579] = f[314] && !f[353] && !f[373] && !f[495];
	assign leaf[9580] = f[314] && !f[353] && !f[373] && f[495];
	assign leaf[9581] = f[314] && !f[353] && f[373] && !f[544];
	assign leaf[9582] = f[314] && !f[353] && f[373] && f[544];
	assign leaf[9583] = f[314] && f[353] && !f[681] && !f[433];
	assign leaf[9584] = f[314] && f[353] && !f[681] && f[433];
	assign leaf[9585] = f[314] && f[353] && f[681];
	
	// Tree 689, Classifier 9, Iteration: 68
	assign leaf[9586] = !f[323] && !f[401] && !f[427] && !f[375];
	assign leaf[9587] = !f[323] && !f[401] && !f[427] && f[375];
	assign leaf[9588] = !f[323] && !f[401] && f[427] && !f[497];
	assign leaf[9589] = !f[323] && !f[401] && f[427] && f[497];
	assign leaf[9590] = !f[323] && f[401] && !f[717] && !f[348];
	assign leaf[9591] = !f[323] && f[401] && !f[717] && f[348];
	assign leaf[9592] = !f[323] && f[401] && f[717] && !f[237];
	assign leaf[9593] = !f[323] && f[401] && f[717] && f[237];
	assign leaf[9594] = f[323] && !f[298] && !f[185] && !f[239];
	assign leaf[9595] = f[323] && !f[298] && !f[185] && f[239];
	assign leaf[9596] = f[323] && !f[298] && f[185] && !f[240];
	assign leaf[9597] = f[323] && !f[298] && f[185] && f[240];
	assign leaf[9598] = f[323] && f[298] && !f[245] && !f[209];
	assign leaf[9599] = f[323] && f[298] && !f[245] && f[209];
	assign leaf[9600] = f[323] && f[298] && f[245] && !f[405];
	assign leaf[9601] = f[323] && f[298] && f[245] && f[405];
	
	// Tree 690, Classifier 0, Iteration: 69
	assign leaf[9602] = !f[633] && !f[580] && !f[378] && !f[599];
	assign leaf[9603] = !f[633] && !f[580] && !f[378] && f[599];
	assign leaf[9604] = !f[633] && !f[580] && f[378] && !f[435];
	assign leaf[9605] = !f[633] && !f[580] && f[378] && f[435];
	assign leaf[9606] = !f[633] && f[580] && !f[568] && !f[471];
	assign leaf[9607] = !f[633] && f[580] && !f[568] && f[471];
	assign leaf[9608] = !f[633] && f[580] && f[568] && !f[182];
	assign leaf[9609] = !f[633] && f[580] && f[568] && f[182];
	assign leaf[9610] = f[633] && !f[234] && !f[205] && !f[686];
	assign leaf[9611] = f[633] && !f[234] && !f[205] && f[686];
	assign leaf[9612] = f[633] && !f[234] && f[205];
	assign leaf[9613] = f[633] && f[234] && !f[629] && !f[179];
	assign leaf[9614] = f[633] && f[234] && !f[629] && f[179];
	assign leaf[9615] = f[633] && f[234] && f[629] && !f[655];
	assign leaf[9616] = f[633] && f[234] && f[629] && f[655];
	
	// Tree 691, Classifier 1, Iteration: 69
	assign leaf[9617] = !f[102] && !f[213] && !f[269] && !f[321];
	assign leaf[9618] = !f[102] && !f[213] && !f[269] && f[321];
	assign leaf[9619] = !f[102] && !f[213] && f[269] && !f[188];
	assign leaf[9620] = !f[102] && !f[213] && f[269] && f[188];
	assign leaf[9621] = !f[102] && f[213] && !f[296] && !f[129];
	assign leaf[9622] = !f[102] && f[213] && !f[296] && f[129];
	assign leaf[9623] = !f[102] && f[213] && f[296] && !f[152];
	assign leaf[9624] = !f[102] && f[213] && f[296] && f[152];
	assign leaf[9625] = f[102] && !f[213];
	assign leaf[9626] = f[102] && f[213];
	
	// Tree 692, Classifier 2, Iteration: 69
	assign leaf[9627] = !f[570] && !f[480] && !f[525] && !f[415];
	assign leaf[9628] = !f[570] && !f[480] && !f[525] && f[415];
	assign leaf[9629] = !f[570] && !f[480] && f[525] && !f[607];
	assign leaf[9630] = !f[570] && !f[480] && f[525] && f[607];
	assign leaf[9631] = !f[570] && f[480] && !f[459];
	assign leaf[9632] = !f[570] && f[480] && f[459] && !f[440];
	assign leaf[9633] = !f[570] && f[480] && f[459] && f[440];
	assign leaf[9634] = f[570] && !f[453] && !f[485] && !f[568];
	assign leaf[9635] = f[570] && !f[453] && !f[485] && f[568];
	assign leaf[9636] = f[570] && !f[453] && f[485] && !f[400];
	assign leaf[9637] = f[570] && !f[453] && f[485] && f[400];
	assign leaf[9638] = f[570] && f[453] && !f[401] && !f[457];
	assign leaf[9639] = f[570] && f[453] && !f[401] && f[457];
	assign leaf[9640] = f[570] && f[453] && f[401] && !f[319];
	assign leaf[9641] = f[570] && f[453] && f[401] && f[319];
	
	// Tree 693, Classifier 3, Iteration: 69
	assign leaf[9642] = !f[434] && !f[321] && !f[96] && !f[351];
	assign leaf[9643] = !f[434] && !f[321] && !f[96] && f[351];
	assign leaf[9644] = !f[434] && !f[321] && f[96] && !f[549];
	assign leaf[9645] = !f[434] && !f[321] && f[96] && f[549];
	assign leaf[9646] = !f[434] && f[321] && !f[347] && !f[436];
	assign leaf[9647] = !f[434] && f[321] && !f[347] && f[436];
	assign leaf[9648] = !f[434] && f[321] && f[347] && !f[288];
	assign leaf[9649] = !f[434] && f[321] && f[347] && f[288];
	assign leaf[9650] = f[434] && !f[208] && !f[461] && !f[406];
	assign leaf[9651] = f[434] && !f[208] && !f[461] && f[406];
	assign leaf[9652] = f[434] && !f[208] && f[461] && !f[606];
	assign leaf[9653] = f[434] && !f[208] && f[461] && f[606];
	assign leaf[9654] = f[434] && f[208] && !f[572] && !f[516];
	assign leaf[9655] = f[434] && f[208] && !f[572] && f[516];
	assign leaf[9656] = f[434] && f[208] && f[572] && !f[489];
	assign leaf[9657] = f[434] && f[208] && f[572] && f[489];
	
	// Tree 694, Classifier 4, Iteration: 69
	assign leaf[9658] = !f[739] && !f[72] && !f[96] && !f[519];
	assign leaf[9659] = !f[739] && !f[72] && !f[96] && f[519];
	assign leaf[9660] = !f[739] && !f[72] && f[96];
	assign leaf[9661] = !f[739] && f[72];
	assign leaf[9662] = f[739] && !f[438];
	assign leaf[9663] = f[739] && f[438];
	
	// Tree 695, Classifier 5, Iteration: 69
	assign leaf[9664] = !f[465] && !f[409] && !f[379] && !f[496];
	assign leaf[9665] = !f[465] && !f[409] && !f[379] && f[496];
	assign leaf[9666] = !f[465] && !f[409] && f[379] && !f[433];
	assign leaf[9667] = !f[465] && !f[409] && f[379] && f[433];
	assign leaf[9668] = !f[465] && f[409] && !f[294] && !f[579];
	assign leaf[9669] = !f[465] && f[409] && !f[294] && f[579];
	assign leaf[9670] = !f[465] && f[409] && f[294] && !f[298];
	assign leaf[9671] = !f[465] && f[409] && f[294] && f[298];
	assign leaf[9672] = f[465] && !f[355] && !f[296] && !f[376];
	assign leaf[9673] = f[465] && !f[355] && !f[296] && f[376];
	assign leaf[9674] = f[465] && !f[355] && f[296] && !f[301];
	assign leaf[9675] = f[465] && !f[355] && f[296] && f[301];
	assign leaf[9676] = f[465] && f[355] && !f[509] && !f[624];
	assign leaf[9677] = f[465] && f[355] && !f[509] && f[624];
	assign leaf[9678] = f[465] && f[355] && f[509] && !f[190];
	assign leaf[9679] = f[465] && f[355] && f[509] && f[190];
	
	// Tree 696, Classifier 6, Iteration: 69
	assign leaf[9680] = !f[601] && !f[208] && !f[523] && !f[542];
	assign leaf[9681] = !f[601] && !f[208] && !f[523] && f[542];
	assign leaf[9682] = !f[601] && !f[208] && f[523] && !f[263];
	assign leaf[9683] = !f[601] && !f[208] && f[523] && f[263];
	assign leaf[9684] = !f[601] && f[208] && !f[180];
	assign leaf[9685] = !f[601] && f[208] && f[180] && !f[263];
	assign leaf[9686] = !f[601] && f[208] && f[180] && f[263];
	assign leaf[9687] = f[601] && !f[627] && !f[178] && !f[516];
	assign leaf[9688] = f[601] && !f[627] && !f[178] && f[516];
	assign leaf[9689] = f[601] && !f[627] && f[178] && !f[631];
	assign leaf[9690] = f[601] && !f[627] && f[178] && f[631];
	assign leaf[9691] = f[601] && f[627] && !f[127] && !f[209];
	assign leaf[9692] = f[601] && f[627] && !f[127] && f[209];
	assign leaf[9693] = f[601] && f[627] && f[127] && !f[455];
	assign leaf[9694] = f[601] && f[627] && f[127] && f[455];
	
	// Tree 697, Classifier 7, Iteration: 69
	assign leaf[9695] = !f[269] && !f[519] && !f[210] && !f[318];
	assign leaf[9696] = !f[269] && !f[519] && !f[210] && f[318];
	assign leaf[9697] = !f[269] && !f[519] && f[210] && !f[373];
	assign leaf[9698] = !f[269] && !f[519] && f[210] && f[373];
	assign leaf[9699] = !f[269] && f[519] && !f[205] && !f[324];
	assign leaf[9700] = !f[269] && f[519] && !f[205] && f[324];
	assign leaf[9701] = !f[269] && f[519] && f[205] && !f[211];
	assign leaf[9702] = !f[269] && f[519] && f[205] && f[211];
	assign leaf[9703] = f[269] && !f[173] && !f[349] && !f[370];
	assign leaf[9704] = f[269] && !f[173] && !f[349] && f[370];
	assign leaf[9705] = f[269] && !f[173] && f[349] && !f[266];
	assign leaf[9706] = f[269] && !f[173] && f[349] && f[266];
	assign leaf[9707] = f[269] && f[173] && !f[550];
	assign leaf[9708] = f[269] && f[173] && f[550];
	
	// Tree 698, Classifier 8, Iteration: 69
	assign leaf[9709] = !f[627] && !f[634] && !f[682] && !f[572];
	assign leaf[9710] = !f[627] && !f[634] && !f[682] && f[572];
	assign leaf[9711] = !f[627] && !f[634] && f[682] && !f[521];
	assign leaf[9712] = !f[627] && !f[634] && f[682] && f[521];
	assign leaf[9713] = !f[627] && f[634] && !f[574] && !f[601];
	assign leaf[9714] = !f[627] && f[634] && !f[574] && f[601];
	assign leaf[9715] = !f[627] && f[634] && f[574] && !f[512];
	assign leaf[9716] = !f[627] && f[634] && f[574] && f[512];
	assign leaf[9717] = f[627] && !f[654] && !f[635] && !f[687];
	assign leaf[9718] = f[627] && !f[654] && !f[635] && f[687];
	assign leaf[9719] = f[627] && !f[654] && f[635] && !f[207];
	assign leaf[9720] = f[627] && !f[654] && f[635] && f[207];
	assign leaf[9721] = f[627] && f[654] && !f[600] && !f[293];
	assign leaf[9722] = f[627] && f[654] && !f[600] && f[293];
	assign leaf[9723] = f[627] && f[654] && f[600] && !f[623];
	assign leaf[9724] = f[627] && f[654] && f[600] && f[623];
	
	// Tree 699, Classifier 9, Iteration: 69
	assign leaf[9725] = !f[500] && !f[350] && !f[438] && !f[522];
	assign leaf[9726] = !f[500] && !f[350] && !f[438] && f[522];
	assign leaf[9727] = !f[500] && !f[350] && f[438] && !f[493];
	assign leaf[9728] = !f[500] && !f[350] && f[438] && f[493];
	assign leaf[9729] = !f[500] && f[350] && !f[460] && !f[241];
	assign leaf[9730] = !f[500] && f[350] && !f[460] && f[241];
	assign leaf[9731] = !f[500] && f[350] && f[460] && !f[372];
	assign leaf[9732] = !f[500] && f[350] && f[460] && f[372];
	assign leaf[9733] = f[500];
	
	// Tree 700, Classifier 0, Iteration: 70
	assign leaf[9734] = !f[380] && !f[456] && !f[424] && !f[267];
	assign leaf[9735] = !f[380] && !f[456] && !f[424] && f[267];
	assign leaf[9736] = !f[380] && !f[456] && f[424] && !f[439];
	assign leaf[9737] = !f[380] && !f[456] && f[424] && f[439];
	assign leaf[9738] = !f[380] && f[456] && !f[654] && !f[575];
	assign leaf[9739] = !f[380] && f[456] && !f[654] && f[575];
	assign leaf[9740] = !f[380] && f[456] && f[654] && !f[512];
	assign leaf[9741] = !f[380] && f[456] && f[654] && f[512];
	assign leaf[9742] = f[380] && !f[350] && !f[324] && !f[407];
	assign leaf[9743] = f[380] && !f[350] && !f[324] && f[407];
	assign leaf[9744] = f[380] && !f[350] && f[324] && !f[262];
	assign leaf[9745] = f[380] && !f[350] && f[324] && f[262];
	assign leaf[9746] = f[380] && f[350] && !f[154] && !f[512];
	assign leaf[9747] = f[380] && f[350] && !f[154] && f[512];
	assign leaf[9748] = f[380] && f[350] && f[154] && !f[382];
	assign leaf[9749] = f[380] && f[350] && f[154] && f[382];
	
	// Tree 701, Classifier 1, Iteration: 70
	assign leaf[9750] = !f[440] && !f[609] && !f[260] && !f[600];
	assign leaf[9751] = !f[440] && !f[609] && !f[260] && f[600];
	assign leaf[9752] = !f[440] && !f[609] && f[260] && !f[153];
	assign leaf[9753] = !f[440] && !f[609] && f[260] && f[153];
	assign leaf[9754] = !f[440] && f[609] && !f[433] && !f[157];
	assign leaf[9755] = !f[440] && f[609] && !f[433] && f[157];
	assign leaf[9756] = !f[440] && f[609] && f[433] && !f[376];
	assign leaf[9757] = !f[440] && f[609] && f[433] && f[376];
	assign leaf[9758] = f[440];
	
	// Tree 702, Classifier 2, Iteration: 70
	assign leaf[9759] = !f[104] && !f[546] && !f[602] && !f[101];
	assign leaf[9760] = !f[104] && !f[546] && !f[602] && f[101];
	assign leaf[9761] = !f[104] && !f[546] && f[602] && !f[492];
	assign leaf[9762] = !f[104] && !f[546] && f[602] && f[492];
	assign leaf[9763] = !f[104] && f[546] && !f[216] && !f[102];
	assign leaf[9764] = !f[104] && f[546] && !f[216] && f[102];
	assign leaf[9765] = !f[104] && f[546] && f[216] && !f[352];
	assign leaf[9766] = !f[104] && f[546] && f[216] && f[352];
	assign leaf[9767] = f[104] && !f[432];
	assign leaf[9768] = f[104] && f[432];
	
	// Tree 703, Classifier 3, Iteration: 70
	assign leaf[9769] = !f[402] && !f[709] && !f[266] && !f[378];
	assign leaf[9770] = !f[402] && !f[709] && !f[266] && f[378];
	assign leaf[9771] = !f[402] && !f[709] && f[266] && !f[160];
	assign leaf[9772] = !f[402] && !f[709] && f[266] && f[160];
	assign leaf[9773] = !f[402] && f[709] && !f[320] && !f[630];
	assign leaf[9774] = !f[402] && f[709] && !f[320] && f[630];
	assign leaf[9775] = !f[402] && f[709] && f[320];
	assign leaf[9776] = f[402] && !f[512] && !f[482] && !f[349];
	assign leaf[9777] = f[402] && !f[512] && !f[482] && f[349];
	assign leaf[9778] = f[402] && !f[512] && f[482] && !f[434];
	assign leaf[9779] = f[402] && !f[512] && f[482] && f[434];
	assign leaf[9780] = f[402] && f[512] && !f[457] && !f[269];
	assign leaf[9781] = f[402] && f[512] && !f[457] && f[269];
	assign leaf[9782] = f[402] && f[512] && f[457] && !f[454];
	assign leaf[9783] = f[402] && f[512] && f[457] && f[454];
	
	// Tree 704, Classifier 4, Iteration: 70
	assign leaf[9784] = !f[399] && !f[286] && !f[184] && !f[267];
	assign leaf[9785] = !f[399] && !f[286] && !f[184] && f[267];
	assign leaf[9786] = !f[399] && !f[286] && f[184] && !f[214];
	assign leaf[9787] = !f[399] && !f[286] && f[184] && f[214];
	assign leaf[9788] = !f[399] && f[286] && !f[426] && !f[211];
	assign leaf[9789] = !f[399] && f[286] && !f[426] && f[211];
	assign leaf[9790] = !f[399] && f[286] && f[426];
	assign leaf[9791] = f[399] && !f[514] && !f[463] && !f[382];
	assign leaf[9792] = f[399] && !f[514] && !f[463] && f[382];
	assign leaf[9793] = f[399] && !f[514] && f[463] && !f[233];
	assign leaf[9794] = f[399] && !f[514] && f[463] && f[233];
	assign leaf[9795] = f[399] && f[514] && !f[467] && !f[327];
	assign leaf[9796] = f[399] && f[514] && !f[467] && f[327];
	assign leaf[9797] = f[399] && f[514] && f[467] && !f[382];
	assign leaf[9798] = f[399] && f[514] && f[467] && f[382];
	
	// Tree 705, Classifier 5, Iteration: 70
	assign leaf[9799] = !f[120] && !f[630] && !f[714] && !f[270];
	assign leaf[9800] = !f[120] && !f[630] && !f[714] && f[270];
	assign leaf[9801] = !f[120] && !f[630] && f[714] && !f[296];
	assign leaf[9802] = !f[120] && !f[630] && f[714] && f[296];
	assign leaf[9803] = !f[120] && f[630] && !f[483] && !f[628];
	assign leaf[9804] = !f[120] && f[630] && !f[483] && f[628];
	assign leaf[9805] = !f[120] && f[630] && f[483] && !f[345];
	assign leaf[9806] = !f[120] && f[630] && f[483] && f[345];
	assign leaf[9807] = f[120] && !f[231] && !f[553];
	assign leaf[9808] = f[120] && !f[231] && f[553];
	assign leaf[9809] = f[120] && f[231];
	
	// Tree 706, Classifier 6, Iteration: 70
	assign leaf[9810] = !f[236] && !f[181] && !f[656] && !f[480];
	assign leaf[9811] = !f[236] && !f[181] && !f[656] && f[480];
	assign leaf[9812] = !f[236] && !f[181] && f[656] && !f[547];
	assign leaf[9813] = !f[236] && !f[181] && f[656] && f[547];
	assign leaf[9814] = !f[236] && f[181] && !f[516] && !f[357];
	assign leaf[9815] = !f[236] && f[181] && !f[516] && f[357];
	assign leaf[9816] = !f[236] && f[181] && f[516] && !f[184];
	assign leaf[9817] = !f[236] && f[181] && f[516] && f[184];
	assign leaf[9818] = f[236] && !f[541] && !f[347] && !f[539];
	assign leaf[9819] = f[236] && !f[541] && !f[347] && f[539];
	assign leaf[9820] = f[236] && !f[541] && f[347] && !f[487];
	assign leaf[9821] = f[236] && !f[541] && f[347] && f[487];
	assign leaf[9822] = f[236] && f[541] && !f[401] && !f[371];
	assign leaf[9823] = f[236] && f[541] && !f[401] && f[371];
	assign leaf[9824] = f[236] && f[541] && f[401] && !f[128];
	assign leaf[9825] = f[236] && f[541] && f[401] && f[128];
	
	// Tree 707, Classifier 7, Iteration: 70
	assign leaf[9826] = !f[214] && !f[543] && !f[457] && !f[370];
	assign leaf[9827] = !f[214] && !f[543] && !f[457] && f[370];
	assign leaf[9828] = !f[214] && !f[543] && f[457] && !f[488];
	assign leaf[9829] = !f[214] && !f[543] && f[457] && f[488];
	assign leaf[9830] = !f[214] && f[543] && !f[679] && !f[528];
	assign leaf[9831] = !f[214] && f[543] && !f[679] && f[528];
	assign leaf[9832] = !f[214] && f[543] && f[679];
	assign leaf[9833] = f[214] && !f[577] && !f[269] && !f[323];
	assign leaf[9834] = f[214] && !f[577] && !f[269] && f[323];
	assign leaf[9835] = f[214] && !f[577] && f[269] && !f[236];
	assign leaf[9836] = f[214] && !f[577] && f[269] && f[236];
	assign leaf[9837] = f[214] && f[577] && !f[716] && !f[715];
	assign leaf[9838] = f[214] && f[577] && !f[716] && f[715];
	assign leaf[9839] = f[214] && f[577] && f[716] && !f[261];
	assign leaf[9840] = f[214] && f[577] && f[716] && f[261];
	
	// Tree 708, Classifier 8, Iteration: 70
	assign leaf[9841] = !f[682] && !f[627] && !f[633] && !f[689];
	assign leaf[9842] = !f[682] && !f[627] && !f[633] && f[689];
	assign leaf[9843] = !f[682] && !f[627] && f[633] && !f[513];
	assign leaf[9844] = !f[682] && !f[627] && f[633] && f[513];
	assign leaf[9845] = !f[682] && f[627] && !f[632] && !f[572];
	assign leaf[9846] = !f[682] && f[627] && !f[632] && f[572];
	assign leaf[9847] = !f[682] && f[627] && f[632] && !f[601];
	assign leaf[9848] = !f[682] && f[627] && f[632] && f[601];
	assign leaf[9849] = f[682] && !f[542] && !f[539] && !f[540];
	assign leaf[9850] = f[682] && !f[542] && !f[539] && f[540];
	assign leaf[9851] = f[682] && !f[542] && f[539] && !f[494];
	assign leaf[9852] = f[682] && !f[542] && f[539] && f[494];
	assign leaf[9853] = f[682] && f[542] && !f[661] && !f[405];
	assign leaf[9854] = f[682] && f[542] && !f[661] && f[405];
	assign leaf[9855] = f[682] && f[542] && f[661] && !f[657];
	assign leaf[9856] = f[682] && f[542] && f[661] && f[657];
	
	// Tree 709, Classifier 9, Iteration: 70
	assign leaf[9857] = !f[734] && !f[247] && !f[122] && !f[228];
	assign leaf[9858] = !f[734] && !f[247] && !f[122] && f[228];
	assign leaf[9859] = !f[734] && !f[247] && f[122];
	assign leaf[9860] = !f[734] && f[247] && !f[215] && !f[514];
	assign leaf[9861] = !f[734] && f[247] && !f[215] && f[514];
	assign leaf[9862] = !f[734] && f[247] && f[215] && !f[404];
	assign leaf[9863] = !f[734] && f[247] && f[215] && f[404];
	assign leaf[9864] = f[734] && !f[624];
	assign leaf[9865] = f[734] && f[624];
	
	// Tree 710, Classifier 0, Iteration: 71
	assign leaf[9866] = !f[688] && !f[152] && !f[654] && !f[275];
	assign leaf[9867] = !f[688] && !f[152] && !f[654] && f[275];
	assign leaf[9868] = !f[688] && !f[152] && f[654] && !f[157];
	assign leaf[9869] = !f[688] && !f[152] && f[654] && f[157];
	assign leaf[9870] = !f[688] && f[152] && !f[349] && !f[293];
	assign leaf[9871] = !f[688] && f[152] && !f[349] && f[293];
	assign leaf[9872] = !f[688] && f[152] && f[349] && !f[238];
	assign leaf[9873] = !f[688] && f[152] && f[349] && f[238];
	assign leaf[9874] = f[688] && !f[657];
	assign leaf[9875] = f[688] && f[657] && !f[231];
	assign leaf[9876] = f[688] && f[657] && f[231];
	
	// Tree 711, Classifier 1, Iteration: 71
	assign leaf[9877] = !f[606] && !f[289] && !f[151] && !f[99];
	assign leaf[9878] = !f[606] && !f[289] && !f[151] && f[99];
	assign leaf[9879] = !f[606] && !f[289] && f[151] && !f[236];
	assign leaf[9880] = !f[606] && !f[289] && f[151] && f[236];
	assign leaf[9881] = !f[606] && f[289];
	assign leaf[9882] = f[606] && !f[491] && !f[379] && !f[461];
	assign leaf[9883] = f[606] && !f[491] && !f[379] && f[461];
	assign leaf[9884] = f[606] && !f[491] && f[379] && !f[626];
	assign leaf[9885] = f[606] && !f[491] && f[379] && f[626];
	assign leaf[9886] = f[606] && f[491] && !f[373] && !f[576];
	assign leaf[9887] = f[606] && f[491] && !f[373] && f[576];
	assign leaf[9888] = f[606] && f[491] && f[373];
	
	// Tree 712, Classifier 2, Iteration: 71
	assign leaf[9889] = !f[276] && !f[378] && !f[400] && !f[275];
	assign leaf[9890] = !f[276] && !f[378] && !f[400] && f[275];
	assign leaf[9891] = !f[276] && !f[378] && f[400] && !f[404];
	assign leaf[9892] = !f[276] && !f[378] && f[400] && f[404];
	assign leaf[9893] = !f[276] && f[378] && !f[214] && !f[658];
	assign leaf[9894] = !f[276] && f[378] && !f[214] && f[658];
	assign leaf[9895] = !f[276] && f[378] && f[214] && !f[100];
	assign leaf[9896] = !f[276] && f[378] && f[214] && f[100];
	assign leaf[9897] = f[276];
	
	// Tree 713, Classifier 3, Iteration: 71
	assign leaf[9898] = !f[712] && !f[718] && !f[626] && !f[683];
	assign leaf[9899] = !f[712] && !f[718] && !f[626] && f[683];
	assign leaf[9900] = !f[712] && !f[718] && f[626] && !f[426];
	assign leaf[9901] = !f[712] && !f[718] && f[626] && f[426];
	assign leaf[9902] = !f[712] && f[718] && !f[489] && !f[459];
	assign leaf[9903] = !f[712] && f[718] && !f[489] && f[459];
	assign leaf[9904] = !f[712] && f[718] && f[489] && !f[493];
	assign leaf[9905] = !f[712] && f[718] && f[489] && f[493];
	assign leaf[9906] = f[712] && !f[375] && !f[409] && !f[433];
	assign leaf[9907] = f[712] && !f[375] && !f[409] && f[433];
	assign leaf[9908] = f[712] && !f[375] && f[409] && !f[430];
	assign leaf[9909] = f[712] && !f[375] && f[409] && f[430];
	assign leaf[9910] = f[712] && f[375] && !f[322] && !f[263];
	assign leaf[9911] = f[712] && f[375] && !f[322] && f[263];
	assign leaf[9912] = f[712] && f[375] && f[322] && !f[319];
	assign leaf[9913] = f[712] && f[375] && f[322] && f[319];
	
	// Tree 714, Classifier 4, Iteration: 71
	assign leaf[9914] = !f[738] && !f[741] && !f[184] && !f[240];
	assign leaf[9915] = !f[738] && !f[741] && !f[184] && f[240];
	assign leaf[9916] = !f[738] && !f[741] && f[184] && !f[240];
	assign leaf[9917] = !f[738] && !f[741] && f[184] && f[240];
	assign leaf[9918] = !f[738] && f[741] && !f[264];
	assign leaf[9919] = !f[738] && f[741] && f[264];
	assign leaf[9920] = f[738];
	
	// Tree 715, Classifier 5, Iteration: 71
	assign leaf[9921] = !f[382] && !f[440] && !f[301] && !f[324];
	assign leaf[9922] = !f[382] && !f[440] && !f[301] && f[324];
	assign leaf[9923] = !f[382] && !f[440] && f[301] && !f[186];
	assign leaf[9924] = !f[382] && !f[440] && f[301] && f[186];
	assign leaf[9925] = !f[382] && f[440] && !f[484] && !f[302];
	assign leaf[9926] = !f[382] && f[440] && !f[484] && f[302];
	assign leaf[9927] = !f[382] && f[440] && f[484] && !f[383];
	assign leaf[9928] = !f[382] && f[440] && f[484] && f[383];
	assign leaf[9929] = f[382] && !f[524] && !f[349] && !f[483];
	assign leaf[9930] = f[382] && !f[524] && !f[349] && f[483];
	assign leaf[9931] = f[382] && !f[524] && f[349] && !f[292];
	assign leaf[9932] = f[382] && !f[524] && f[349] && f[292];
	assign leaf[9933] = f[382] && f[524] && !f[490] && !f[233];
	assign leaf[9934] = f[382] && f[524] && !f[490] && f[233];
	assign leaf[9935] = f[382] && f[524] && f[490] && !f[240];
	assign leaf[9936] = f[382] && f[524] && f[490] && f[240];
	
	// Tree 716, Classifier 6, Iteration: 71
	assign leaf[9937] = !f[622] && !f[101] && !f[212] && !f[320];
	assign leaf[9938] = !f[622] && !f[101] && !f[212] && f[320];
	assign leaf[9939] = !f[622] && !f[101] && f[212] && !f[486];
	assign leaf[9940] = !f[622] && !f[101] && f[212] && f[486];
	assign leaf[9941] = !f[622] && f[101] && !f[211] && !f[580];
	assign leaf[9942] = !f[622] && f[101] && !f[211] && f[580];
	assign leaf[9943] = !f[622] && f[101] && f[211] && !f[631];
	assign leaf[9944] = !f[622] && f[101] && f[211] && f[631];
	assign leaf[9945] = f[622];
	
	// Tree 717, Classifier 7, Iteration: 71
	assign leaf[9946] = !f[494] && !f[605] && !f[690] && !f[575];
	assign leaf[9947] = !f[494] && !f[605] && !f[690] && f[575];
	assign leaf[9948] = !f[494] && !f[605] && f[690] && !f[440];
	assign leaf[9949] = !f[494] && !f[605] && f[690] && f[440];
	assign leaf[9950] = !f[494] && f[605] && !f[285] && !f[455];
	assign leaf[9951] = !f[494] && f[605] && !f[285] && f[455];
	assign leaf[9952] = !f[494] && f[605] && f[285] && !f[579];
	assign leaf[9953] = !f[494] && f[605] && f[285] && f[579];
	assign leaf[9954] = f[494] && !f[571] && !f[655] && !f[576];
	assign leaf[9955] = f[494] && !f[571] && !f[655] && f[576];
	assign leaf[9956] = f[494] && !f[571] && f[655] && !f[518];
	assign leaf[9957] = f[494] && !f[571] && f[655] && f[518];
	assign leaf[9958] = f[494] && f[571] && !f[654] && !f[173];
	assign leaf[9959] = f[494] && f[571] && !f[654] && f[173];
	assign leaf[9960] = f[494] && f[571] && f[654] && !f[516];
	assign leaf[9961] = f[494] && f[571] && f[654] && f[516];
	
	// Tree 718, Classifier 8, Iteration: 71
	assign leaf[9962] = !f[542] && !f[512] && !f[653] && !f[545];
	assign leaf[9963] = !f[542] && !f[512] && !f[653] && f[545];
	assign leaf[9964] = !f[542] && !f[512] && f[653] && !f[509];
	assign leaf[9965] = !f[542] && !f[512] && f[653] && f[509];
	assign leaf[9966] = !f[542] && f[512] && !f[379] && !f[635];
	assign leaf[9967] = !f[542] && f[512] && !f[379] && f[635];
	assign leaf[9968] = !f[542] && f[512] && f[379] && !f[604];
	assign leaf[9969] = !f[542] && f[512] && f[379] && f[604];
	assign leaf[9970] = f[542] && !f[512] && !f[324] && !f[576];
	assign leaf[9971] = f[542] && !f[512] && !f[324] && f[576];
	assign leaf[9972] = f[542] && !f[512] && f[324] && !f[241];
	assign leaf[9973] = f[542] && !f[512] && f[324] && f[241];
	assign leaf[9974] = f[542] && f[512] && !f[458] && !f[576];
	assign leaf[9975] = f[542] && f[512] && !f[458] && f[576];
	assign leaf[9976] = f[542] && f[512] && f[458] && !f[682];
	assign leaf[9977] = f[542] && f[512] && f[458] && f[682];
	
	// Tree 719, Classifier 9, Iteration: 71
	assign leaf[9978] = !f[566] && !f[175] && !f[639] && !f[524];
	assign leaf[9979] = !f[566] && !f[175] && !f[639] && f[524];
	assign leaf[9980] = !f[566] && !f[175] && f[639] && !f[426];
	assign leaf[9981] = !f[566] && !f[175] && f[639] && f[426];
	assign leaf[9982] = !f[566] && f[175] && !f[690];
	assign leaf[9983] = !f[566] && f[175] && f[690];
	assign leaf[9984] = f[566] && !f[551];
	assign leaf[9985] = f[566] && f[551] && !f[320] && !f[315];
	assign leaf[9986] = f[566] && f[551] && !f[320] && f[315];
	assign leaf[9987] = f[566] && f[551] && f[320];
	
	// Tree 720, Classifier 0, Iteration: 72
	assign leaf[9988] = !f[466] && !f[213] && !f[293] && !f[517];
	assign leaf[9989] = !f[466] && !f[213] && !f[293] && f[517];
	assign leaf[9990] = !f[466] && !f[213] && f[293] && !f[521];
	assign leaf[9991] = !f[466] && !f[213] && f[293] && f[521];
	assign leaf[9992] = !f[466] && f[213] && !f[513] && !f[410];
	assign leaf[9993] = !f[466] && f[213] && !f[513] && f[410];
	assign leaf[9994] = !f[466] && f[213] && f[513] && !f[524];
	assign leaf[9995] = !f[466] && f[213] && f[513] && f[524];
	assign leaf[9996] = f[466] && !f[688] && !f[379] && !f[551];
	assign leaf[9997] = f[466] && !f[688] && !f[379] && f[551];
	assign leaf[9998] = f[466] && !f[688] && f[379] && !f[659];
	assign leaf[9999] = f[466] && !f[688] && f[379] && f[659];
	assign leaf[10000] = f[466] && f[688];
	
	// Tree 721, Classifier 1, Iteration: 72
	assign leaf[10001] = !f[578] && !f[177] && !f[658] && !f[601];
	assign leaf[10002] = !f[578] && !f[177] && !f[658] && f[601];
	assign leaf[10003] = !f[578] && !f[177] && f[658] && !f[266];
	assign leaf[10004] = !f[578] && !f[177] && f[658] && f[266];
	assign leaf[10005] = !f[578] && f[177] && !f[605];
	assign leaf[10006] = !f[578] && f[177] && f[605];
	assign leaf[10007] = f[578] && !f[515] && !f[576] && !f[182];
	assign leaf[10008] = f[578] && !f[515] && !f[576] && f[182];
	assign leaf[10009] = f[578] && !f[515] && f[576] && !f[317];
	assign leaf[10010] = f[578] && !f[515] && f[576] && f[317];
	assign leaf[10011] = f[578] && f[515] && !f[540] && !f[375];
	assign leaf[10012] = f[578] && f[515] && !f[540] && f[375];
	assign leaf[10013] = f[578] && f[515] && f[540];
	
	// Tree 722, Classifier 2, Iteration: 72
	assign leaf[10014] = !f[712] && !f[677] && !f[322] && !f[657];
	assign leaf[10015] = !f[712] && !f[677] && !f[322] && f[657];
	assign leaf[10016] = !f[712] && !f[677] && f[322] && !f[325];
	assign leaf[10017] = !f[712] && !f[677] && f[322] && f[325];
	assign leaf[10018] = !f[712] && f[677];
	assign leaf[10019] = f[712] && !f[406];
	assign leaf[10020] = f[712] && f[406];
	
	// Tree 723, Classifier 3, Iteration: 72
	assign leaf[10021] = !f[373] && !f[689] && !f[740] && !f[715];
	assign leaf[10022] = !f[373] && !f[689] && !f[740] && f[715];
	assign leaf[10023] = !f[373] && !f[689] && f[740];
	assign leaf[10024] = !f[373] && f[689] && !f[575] && !f[519];
	assign leaf[10025] = !f[373] && f[689] && !f[575] && f[519];
	assign leaf[10026] = !f[373] && f[689] && f[575] && !f[492];
	assign leaf[10027] = !f[373] && f[689] && f[575] && f[492];
	assign leaf[10028] = f[373] && !f[320] && !f[264] && !f[233];
	assign leaf[10029] = f[373] && !f[320] && !f[264] && f[233];
	assign leaf[10030] = f[373] && !f[320] && f[264] && !f[239];
	assign leaf[10031] = f[373] && !f[320] && f[264] && f[239];
	assign leaf[10032] = f[373] && f[320] && !f[298] && !f[216];
	assign leaf[10033] = f[373] && f[320] && !f[298] && f[216];
	assign leaf[10034] = f[373] && f[320] && f[298] && !f[155];
	assign leaf[10035] = f[373] && f[320] && f[298] && f[155];
	
	// Tree 724, Classifier 4, Iteration: 72
	assign leaf[10036] = !f[179] && !f[153] && !f[178] && !f[263];
	assign leaf[10037] = !f[179] && !f[153] && !f[178] && f[263];
	assign leaf[10038] = !f[179] && !f[153] && f[178] && !f[269];
	assign leaf[10039] = !f[179] && !f[153] && f[178] && f[269];
	assign leaf[10040] = !f[179] && f[153] && !f[551] && !f[464];
	assign leaf[10041] = !f[179] && f[153] && !f[551] && f[464];
	assign leaf[10042] = !f[179] && f[153] && f[551] && !f[520];
	assign leaf[10043] = !f[179] && f[153] && f[551] && f[520];
	assign leaf[10044] = f[179] && !f[155] && !f[204] && !f[213];
	assign leaf[10045] = f[179] && !f[155] && !f[204] && f[213];
	assign leaf[10046] = f[179] && !f[155] && f[204] && !f[436];
	assign leaf[10047] = f[179] && !f[155] && f[204] && f[436];
	assign leaf[10048] = f[179] && f[155] && !f[540] && !f[267];
	assign leaf[10049] = f[179] && f[155] && !f[540] && f[267];
	assign leaf[10050] = f[179] && f[155] && f[540];
	
	// Tree 725, Classifier 5, Iteration: 72
	assign leaf[10051] = !f[102] && !f[584] && !f[483] && !f[625];
	assign leaf[10052] = !f[102] && !f[584] && !f[483] && f[625];
	assign leaf[10053] = !f[102] && !f[584] && f[483] && !f[428];
	assign leaf[10054] = !f[102] && !f[584] && f[483] && f[428];
	assign leaf[10055] = !f[102] && f[584] && !f[290];
	assign leaf[10056] = !f[102] && f[584] && f[290];
	assign leaf[10057] = f[102] && !f[603];
	assign leaf[10058] = f[102] && f[603] && !f[401] && !f[431];
	assign leaf[10059] = f[102] && f[603] && !f[401] && f[431];
	assign leaf[10060] = f[102] && f[603] && f[401] && !f[237];
	assign leaf[10061] = f[102] && f[603] && f[401] && f[237];
	
	// Tree 726, Classifier 6, Iteration: 72
	assign leaf[10062] = !f[269] && !f[301] && !f[232] && !f[399];
	assign leaf[10063] = !f[269] && !f[301] && !f[232] && f[399];
	assign leaf[10064] = !f[269] && !f[301] && f[232] && !f[347];
	assign leaf[10065] = !f[269] && !f[301] && f[232] && f[347];
	assign leaf[10066] = !f[269] && f[301] && !f[299] && !f[359];
	assign leaf[10067] = !f[269] && f[301] && !f[299] && f[359];
	assign leaf[10068] = !f[269] && f[301] && f[299] && !f[383];
	assign leaf[10069] = !f[269] && f[301] && f[299] && f[383];
	assign leaf[10070] = f[269] && !f[662] && !f[164] && !f[604];
	assign leaf[10071] = f[269] && !f[662] && !f[164] && f[604];
	assign leaf[10072] = f[269] && !f[662] && f[164] && !f[319];
	assign leaf[10073] = f[269] && !f[662] && f[164] && f[319];
	assign leaf[10074] = f[269] && f[662];
	
	// Tree 727, Classifier 7, Iteration: 72
	assign leaf[10075] = !f[359] && !f[663] && !f[320] && !f[317];
	assign leaf[10076] = !f[359] && !f[663] && !f[320] && f[317];
	assign leaf[10077] = !f[359] && !f[663] && f[320] && !f[318];
	assign leaf[10078] = !f[359] && !f[663] && f[320] && f[318];
	assign leaf[10079] = !f[359] && f[663] && !f[577] && !f[178];
	assign leaf[10080] = !f[359] && f[663] && !f[577] && f[178];
	assign leaf[10081] = !f[359] && f[663] && f[577] && !f[516];
	assign leaf[10082] = !f[359] && f[663] && f[577] && f[516];
	assign leaf[10083] = f[359] && !f[456] && !f[369];
	assign leaf[10084] = f[359] && !f[456] && f[369];
	assign leaf[10085] = f[359] && f[456] && !f[485];
	assign leaf[10086] = f[359] && f[456] && f[485];
	
	// Tree 728, Classifier 8, Iteration: 72
	assign leaf[10087] = !f[176] && !f[292] && !f[265] && !f[598];
	assign leaf[10088] = !f[176] && !f[292] && !f[265] && f[598];
	assign leaf[10089] = !f[176] && !f[292] && f[265] && !f[239];
	assign leaf[10090] = !f[176] && !f[292] && f[265] && f[239];
	assign leaf[10091] = !f[176] && f[292] && !f[349] && !f[685];
	assign leaf[10092] = !f[176] && f[292] && !f[349] && f[685];
	assign leaf[10093] = !f[176] && f[292] && f[349] && !f[238];
	assign leaf[10094] = !f[176] && f[292] && f[349] && f[238];
	assign leaf[10095] = f[176] && !f[657] && !f[631] && !f[183];
	assign leaf[10096] = f[176] && !f[657] && !f[631] && f[183];
	assign leaf[10097] = f[176] && !f[657] && f[631] && !f[607];
	assign leaf[10098] = f[176] && !f[657] && f[631] && f[607];
	assign leaf[10099] = f[176] && f[657] && !f[321] && !f[630];
	assign leaf[10100] = f[176] && f[657] && !f[321] && f[630];
	assign leaf[10101] = f[176] && f[657] && f[321] && !f[346];
	assign leaf[10102] = f[176] && f[657] && f[321] && f[346];
	
	// Tree 729, Classifier 9, Iteration: 72
	assign leaf[10103] = !f[381] && !f[432] && !f[491] && !f[206];
	assign leaf[10104] = !f[381] && !f[432] && !f[491] && f[206];
	assign leaf[10105] = !f[381] && !f[432] && f[491] && !f[156];
	assign leaf[10106] = !f[381] && !f[432] && f[491] && f[156];
	assign leaf[10107] = !f[381] && f[432] && !f[374] && !f[460];
	assign leaf[10108] = !f[381] && f[432] && !f[374] && f[460];
	assign leaf[10109] = !f[381] && f[432] && f[374] && !f[514];
	assign leaf[10110] = !f[381] && f[432] && f[374] && f[514];
	assign leaf[10111] = f[381] && !f[437] && !f[520] && !f[263];
	assign leaf[10112] = f[381] && !f[437] && !f[520] && f[263];
	assign leaf[10113] = f[381] && !f[437] && f[520] && !f[490];
	assign leaf[10114] = f[381] && !f[437] && f[520] && f[490];
	assign leaf[10115] = f[381] && f[437] && !f[210] && !f[547];
	assign leaf[10116] = f[381] && f[437] && !f[210] && f[547];
	assign leaf[10117] = f[381] && f[437] && f[210] && !f[265];
	assign leaf[10118] = f[381] && f[437] && f[210] && f[265];
	
	// Tree 730, Classifier 0, Iteration: 73
	assign leaf[10119] = !f[683] && !f[714] && !f[183] && !f[609];
	assign leaf[10120] = !f[683] && !f[714] && !f[183] && f[609];
	assign leaf[10121] = !f[683] && !f[714] && f[183] && !f[630];
	assign leaf[10122] = !f[683] && !f[714] && f[183] && f[630];
	assign leaf[10123] = !f[683] && f[714];
	assign leaf[10124] = f[683] && !f[185];
	assign leaf[10125] = f[683] && f[185] && !f[490] && !f[272];
	assign leaf[10126] = f[683] && f[185] && !f[490] && f[272];
	assign leaf[10127] = f[683] && f[185] && f[490];
	
	// Tree 731, Classifier 1, Iteration: 73
	assign leaf[10128] = !f[381] && !f[464] && !f[324] && !f[177];
	assign leaf[10129] = !f[381] && !f[464] && !f[324] && f[177];
	assign leaf[10130] = !f[381] && !f[464] && f[324] && !f[264];
	assign leaf[10131] = !f[381] && !f[464] && f[324] && f[264];
	assign leaf[10132] = !f[381] && f[464] && !f[237] && !f[232];
	assign leaf[10133] = !f[381] && f[464] && !f[237] && f[232];
	assign leaf[10134] = !f[381] && f[464] && f[237] && !f[208];
	assign leaf[10135] = !f[381] && f[464] && f[237] && f[208];
	assign leaf[10136] = f[381] && !f[297] && !f[213] && !f[436];
	assign leaf[10137] = f[381] && !f[297] && !f[213] && f[436];
	assign leaf[10138] = f[381] && !f[297] && f[213] && !f[327];
	assign leaf[10139] = f[381] && !f[297] && f[213] && f[327];
	assign leaf[10140] = f[381] && f[297] && !f[268] && !f[595];
	assign leaf[10141] = f[381] && f[297] && !f[268] && f[595];
	assign leaf[10142] = f[381] && f[297] && f[268] && !f[152];
	assign leaf[10143] = f[381] && f[297] && f[268] && f[152];
	
	// Tree 732, Classifier 2, Iteration: 73
	assign leaf[10144] = !f[219] && !f[514] && !f[460] && !f[715];
	assign leaf[10145] = !f[219] && !f[514] && !f[460] && f[715];
	assign leaf[10146] = !f[219] && !f[514] && f[460] && !f[509];
	assign leaf[10147] = !f[219] && !f[514] && f[460] && f[509];
	assign leaf[10148] = !f[219] && f[514] && !f[259] && !f[293];
	assign leaf[10149] = !f[219] && f[514] && !f[259] && f[293];
	assign leaf[10150] = !f[219] && f[514] && f[259] && !f[455];
	assign leaf[10151] = !f[219] && f[514] && f[259] && f[455];
	assign leaf[10152] = f[219] && !f[622] && !f[599];
	assign leaf[10153] = f[219] && !f[622] && f[599];
	assign leaf[10154] = f[219] && f[622] && !f[603];
	assign leaf[10155] = f[219] && f[622] && f[603];
	
	// Tree 733, Classifier 3, Iteration: 73
	assign leaf[10156] = !f[331] && !f[676] && !f[479] && !f[604];
	assign leaf[10157] = !f[331] && !f[676] && !f[479] && f[604];
	assign leaf[10158] = !f[331] && !f[676] && f[479] && !f[426];
	assign leaf[10159] = !f[331] && !f[676] && f[479] && f[426];
	assign leaf[10160] = !f[331] && f[676];
	assign leaf[10161] = f[331] && !f[234];
	assign leaf[10162] = f[331] && f[234];
	
	// Tree 734, Classifier 4, Iteration: 73
	assign leaf[10163] = !f[637] && !f[444] && !f[570] && !f[624];
	assign leaf[10164] = !f[637] && !f[444] && !f[570] && f[624];
	assign leaf[10165] = !f[637] && !f[444] && f[570] && !f[400];
	assign leaf[10166] = !f[637] && !f[444] && f[570] && f[400];
	assign leaf[10167] = !f[637] && f[444] && !f[298] && !f[211];
	assign leaf[10168] = !f[637] && f[444] && !f[298] && f[211];
	assign leaf[10169] = !f[637] && f[444] && f[298] && !f[454];
	assign leaf[10170] = !f[637] && f[444] && f[298] && f[454];
	assign leaf[10171] = f[637] && !f[234] && !f[522];
	assign leaf[10172] = f[637] && !f[234] && f[522] && !f[399];
	assign leaf[10173] = f[637] && !f[234] && f[522] && f[399];
	assign leaf[10174] = f[637] && f[234] && !f[453] && !f[210];
	assign leaf[10175] = f[637] && f[234] && !f[453] && f[210];
	assign leaf[10176] = f[637] && f[234] && f[453];
	
	// Tree 735, Classifier 5, Iteration: 73
	assign leaf[10177] = !f[145] && !f[285] && !f[380] && !f[353];
	assign leaf[10178] = !f[145] && !f[285] && !f[380] && f[353];
	assign leaf[10179] = !f[145] && !f[285] && f[380] && !f[377];
	assign leaf[10180] = !f[145] && !f[285] && f[380] && f[377];
	assign leaf[10181] = !f[145] && f[285] && !f[371] && !f[185];
	assign leaf[10182] = !f[145] && f[285] && !f[371] && f[185];
	assign leaf[10183] = !f[145] && f[285] && f[371] && !f[527];
	assign leaf[10184] = !f[145] && f[285] && f[371] && f[527];
	assign leaf[10185] = f[145];
	
	// Tree 736, Classifier 6, Iteration: 73
	assign leaf[10186] = !f[432] && !f[214] && !f[349] && !f[155];
	assign leaf[10187] = !f[432] && !f[214] && !f[349] && f[155];
	assign leaf[10188] = !f[432] && !f[214] && f[349] && !f[457];
	assign leaf[10189] = !f[432] && !f[214] && f[349] && f[457];
	assign leaf[10190] = !f[432] && f[214] && !f[238] && !f[433];
	assign leaf[10191] = !f[432] && f[214] && !f[238] && f[433];
	assign leaf[10192] = !f[432] && f[214] && f[238] && !f[159];
	assign leaf[10193] = !f[432] && f[214] && f[238] && f[159];
	assign leaf[10194] = f[432] && !f[516] && !f[541] && !f[510];
	assign leaf[10195] = f[432] && !f[516] && !f[541] && f[510];
	assign leaf[10196] = f[432] && !f[516] && f[541] && !f[326];
	assign leaf[10197] = f[432] && !f[516] && f[541] && f[326];
	assign leaf[10198] = f[432] && f[516] && !f[155] && !f[237];
	assign leaf[10199] = f[432] && f[516] && !f[155] && f[237];
	assign leaf[10200] = f[432] && f[516] && f[155] && !f[244];
	assign leaf[10201] = f[432] && f[516] && f[155] && f[244];
	
	// Tree 737, Classifier 7, Iteration: 73
	assign leaf[10202] = !f[154] && !f[159] && !f[461] && !f[378];
	assign leaf[10203] = !f[154] && !f[159] && !f[461] && f[378];
	assign leaf[10204] = !f[154] && !f[159] && f[461] && !f[378];
	assign leaf[10205] = !f[154] && !f[159] && f[461] && f[378];
	assign leaf[10206] = !f[154] && f[159] && !f[263];
	assign leaf[10207] = !f[154] && f[159] && f[263];
	assign leaf[10208] = f[154] && !f[236] && !f[262] && !f[260];
	assign leaf[10209] = f[154] && !f[236] && !f[262] && f[260];
	assign leaf[10210] = f[154] && !f[236] && f[262];
	assign leaf[10211] = f[154] && f[236] && !f[684] && !f[232];
	assign leaf[10212] = f[154] && f[236] && !f[684] && f[232];
	assign leaf[10213] = f[154] && f[236] && f[684] && !f[234];
	assign leaf[10214] = f[154] && f[236] && f[684] && f[234];
	
	// Tree 738, Classifier 8, Iteration: 73
	assign leaf[10215] = !f[214] && !f[265] && !f[461] && !f[345];
	assign leaf[10216] = !f[214] && !f[265] && !f[461] && f[345];
	assign leaf[10217] = !f[214] && !f[265] && f[461] && !f[320];
	assign leaf[10218] = !f[214] && !f[265] && f[461] && f[320];
	assign leaf[10219] = !f[214] && f[265] && !f[320] && !f[570];
	assign leaf[10220] = !f[214] && f[265] && !f[320] && f[570];
	assign leaf[10221] = !f[214] && f[265] && f[320] && !f[162];
	assign leaf[10222] = !f[214] && f[265] && f[320] && f[162];
	assign leaf[10223] = f[214] && !f[408] && !f[216] && !f[547];
	assign leaf[10224] = f[214] && !f[408] && !f[216] && f[547];
	assign leaf[10225] = f[214] && !f[408] && f[216] && !f[576];
	assign leaf[10226] = f[214] && !f[408] && f[216] && f[576];
	assign leaf[10227] = f[214] && f[408] && !f[603] && !f[491];
	assign leaf[10228] = f[214] && f[408] && !f[603] && f[491];
	assign leaf[10229] = f[214] && f[408] && f[603] && !f[398];
	assign leaf[10230] = f[214] && f[408] && f[603] && f[398];
	
	// Tree 739, Classifier 9, Iteration: 73
	assign leaf[10231] = !f[734] && !f[368] && !f[374] && !f[400];
	assign leaf[10232] = !f[734] && !f[368] && !f[374] && f[400];
	assign leaf[10233] = !f[734] && !f[368] && f[374] && !f[400];
	assign leaf[10234] = !f[734] && !f[368] && f[374] && f[400];
	assign leaf[10235] = !f[734] && f[368] && !f[347] && !f[270];
	assign leaf[10236] = !f[734] && f[368] && !f[347] && f[270];
	assign leaf[10237] = !f[734] && f[368] && f[347];
	assign leaf[10238] = f[734] && !f[321];
	assign leaf[10239] = f[734] && f[321];
	
	// Tree 740, Classifier 0, Iteration: 74
	assign leaf[10240] = !f[427] && !f[597] && !f[571] && !f[317];
	assign leaf[10241] = !f[427] && !f[597] && !f[571] && f[317];
	assign leaf[10242] = !f[427] && !f[597] && f[571] && !f[263];
	assign leaf[10243] = !f[427] && !f[597] && f[571] && f[263];
	assign leaf[10244] = !f[427] && f[597] && !f[516] && !f[324];
	assign leaf[10245] = !f[427] && f[597] && !f[516] && f[324];
	assign leaf[10246] = !f[427] && f[597] && f[516] && !f[406];
	assign leaf[10247] = !f[427] && f[597] && f[516] && f[406];
	assign leaf[10248] = f[427] && !f[569] && !f[431] && !f[324];
	assign leaf[10249] = f[427] && !f[569] && !f[431] && f[324];
	assign leaf[10250] = f[427] && !f[569] && f[431];
	assign leaf[10251] = f[427] && f[569] && !f[458] && !f[548];
	assign leaf[10252] = f[427] && f[569] && !f[458] && f[548];
	assign leaf[10253] = f[427] && f[569] && f[458] && !f[440];
	assign leaf[10254] = f[427] && f[569] && f[458] && f[440];
	
	// Tree 741, Classifier 1, Iteration: 74
	assign leaf[10255] = !f[555] && !f[96] && !f[378] && !f[517];
	assign leaf[10256] = !f[555] && !f[96] && !f[378] && f[517];
	assign leaf[10257] = !f[555] && !f[96] && f[378] && !f[322];
	assign leaf[10258] = !f[555] && !f[96] && f[378] && f[322];
	assign leaf[10259] = !f[555] && f[96];
	assign leaf[10260] = f[555] && !f[568];
	assign leaf[10261] = f[555] && f[568];
	
	// Tree 742, Classifier 2, Iteration: 74
	assign leaf[10262] = !f[411] && !f[173] && !f[356] && !f[463];
	assign leaf[10263] = !f[411] && !f[173] && !f[356] && f[463];
	assign leaf[10264] = !f[411] && !f[173] && f[356] && !f[463];
	assign leaf[10265] = !f[411] && !f[173] && f[356] && f[463];
	assign leaf[10266] = !f[411] && f[173] && !f[258] && !f[544];
	assign leaf[10267] = !f[411] && f[173] && !f[258] && f[544];
	assign leaf[10268] = !f[411] && f[173] && f[258];
	assign leaf[10269] = f[411] && !f[493] && !f[512] && !f[600];
	assign leaf[10270] = f[411] && !f[493] && !f[512] && f[600];
	assign leaf[10271] = f[411] && !f[493] && f[512] && !f[489];
	assign leaf[10272] = f[411] && !f[493] && f[512] && f[489];
	assign leaf[10273] = f[411] && f[493] && !f[518] && !f[148];
	assign leaf[10274] = f[411] && f[493] && !f[518] && f[148];
	assign leaf[10275] = f[411] && f[493] && f[518] && !f[555];
	assign leaf[10276] = f[411] && f[493] && f[518] && f[555];
	
	// Tree 743, Classifier 3, Iteration: 74
	assign leaf[10277] = !f[120] && !f[269] && !f[296] && !f[513];
	assign leaf[10278] = !f[120] && !f[269] && !f[296] && f[513];
	assign leaf[10279] = !f[120] && !f[269] && f[296] && !f[129];
	assign leaf[10280] = !f[120] && !f[269] && f[296] && f[129];
	assign leaf[10281] = !f[120] && f[269] && !f[101] && !f[378];
	assign leaf[10282] = !f[120] && f[269] && !f[101] && f[378];
	assign leaf[10283] = !f[120] && f[269] && f[101] && !f[579];
	assign leaf[10284] = !f[120] && f[269] && f[101] && f[579];
	assign leaf[10285] = f[120] && !f[630];
	assign leaf[10286] = f[120] && f[630] && !f[458] && !f[292];
	assign leaf[10287] = f[120] && f[630] && !f[458] && f[292];
	assign leaf[10288] = f[120] && f[630] && f[458];
	
	// Tree 744, Classifier 4, Iteration: 74
	assign leaf[10289] = !f[601] && !f[657] && !f[441] && !f[459];
	assign leaf[10290] = !f[601] && !f[657] && !f[441] && f[459];
	assign leaf[10291] = !f[601] && !f[657] && f[441] && !f[217];
	assign leaf[10292] = !f[601] && !f[657] && f[441] && f[217];
	assign leaf[10293] = !f[601] && f[657] && !f[437] && !f[267];
	assign leaf[10294] = !f[601] && f[657] && !f[437] && f[267];
	assign leaf[10295] = !f[601] && f[657] && f[437] && !f[547];
	assign leaf[10296] = !f[601] && f[657] && f[437] && f[547];
	assign leaf[10297] = f[601] && !f[518] && !f[399];
	assign leaf[10298] = f[601] && !f[518] && f[399] && !f[240];
	assign leaf[10299] = f[601] && !f[518] && f[399] && f[240];
	assign leaf[10300] = f[601] && f[518] && !f[239] && !f[322];
	assign leaf[10301] = f[601] && f[518] && !f[239] && f[322];
	assign leaf[10302] = f[601] && f[518] && f[239] && !f[468];
	assign leaf[10303] = f[601] && f[518] && f[239] && f[468];
	
	// Tree 745, Classifier 5, Iteration: 74
	assign leaf[10304] = !f[322] && !f[349] && !f[520] && !f[263];
	assign leaf[10305] = !f[322] && !f[349] && !f[520] && f[263];
	assign leaf[10306] = !f[322] && !f[349] && f[520] && !f[490];
	assign leaf[10307] = !f[322] && !f[349] && f[520] && f[490];
	assign leaf[10308] = !f[322] && f[349] && !f[174] && !f[267];
	assign leaf[10309] = !f[322] && f[349] && !f[174] && f[267];
	assign leaf[10310] = !f[322] && f[349] && f[174] && !f[235];
	assign leaf[10311] = !f[322] && f[349] && f[174] && f[235];
	assign leaf[10312] = f[322] && !f[218] && !f[268] && !f[156];
	assign leaf[10313] = f[322] && !f[218] && !f[268] && f[156];
	assign leaf[10314] = f[322] && !f[218] && f[268] && !f[295];
	assign leaf[10315] = f[322] && !f[218] && f[268] && f[295];
	assign leaf[10316] = f[322] && f[218] && !f[160] && !f[273];
	assign leaf[10317] = f[322] && f[218] && !f[160] && f[273];
	assign leaf[10318] = f[322] && f[218] && f[160] && !f[237];
	assign leaf[10319] = f[322] && f[218] && f[160] && f[237];
	
	// Tree 746, Classifier 6, Iteration: 74
	assign leaf[10320] = !f[302] && !f[299] && !f[399] && !f[518];
	assign leaf[10321] = !f[302] && !f[299] && !f[399] && f[518];
	assign leaf[10322] = !f[302] && !f[299] && f[399] && !f[269];
	assign leaf[10323] = !f[302] && !f[299] && f[399] && f[269];
	assign leaf[10324] = !f[302] && f[299] && !f[457] && !f[301];
	assign leaf[10325] = !f[302] && f[299] && !f[457] && f[301];
	assign leaf[10326] = !f[302] && f[299] && f[457] && !f[382];
	assign leaf[10327] = !f[302] && f[299] && f[457] && f[382];
	assign leaf[10328] = f[302] && !f[416] && !f[271] && !f[408];
	assign leaf[10329] = f[302] && !f[416] && !f[271] && f[408];
	assign leaf[10330] = f[302] && !f[416] && f[271] && !f[430];
	assign leaf[10331] = f[302] && !f[416] && f[271] && f[430];
	assign leaf[10332] = f[302] && f[416];
	
	// Tree 747, Classifier 7, Iteration: 74
	assign leaf[10333] = !f[709] && !f[129] && !f[214] && !f[323];
	assign leaf[10334] = !f[709] && !f[129] && !f[214] && f[323];
	assign leaf[10335] = !f[709] && !f[129] && f[214] && !f[320];
	assign leaf[10336] = !f[709] && !f[129] && f[214] && f[320];
	assign leaf[10337] = !f[709] && f[129];
	assign leaf[10338] = f[709] && !f[654] && !f[271];
	assign leaf[10339] = f[709] && !f[654] && f[271];
	assign leaf[10340] = f[709] && f[654] && !f[322] && !f[303];
	assign leaf[10341] = f[709] && f[654] && !f[322] && f[303];
	assign leaf[10342] = f[709] && f[654] && f[322] && !f[329];
	assign leaf[10343] = f[709] && f[654] && f[322] && f[329];
	
	// Tree 748, Classifier 8, Iteration: 74
	assign leaf[10344] = !f[349] && !f[519] && !f[355] && !f[521];
	assign leaf[10345] = !f[349] && !f[519] && !f[355] && f[521];
	assign leaf[10346] = !f[349] && !f[519] && f[355] && !f[326];
	assign leaf[10347] = !f[349] && !f[519] && f[355] && f[326];
	assign leaf[10348] = !f[349] && f[519] && !f[543] && !f[663];
	assign leaf[10349] = !f[349] && f[519] && !f[543] && f[663];
	assign leaf[10350] = !f[349] && f[519] && f[543] && !f[512];
	assign leaf[10351] = !f[349] && f[519] && f[543] && f[512];
	assign leaf[10352] = f[349] && !f[519] && !f[436] && !f[544];
	assign leaf[10353] = f[349] && !f[519] && !f[436] && f[544];
	assign leaf[10354] = f[349] && !f[519] && f[436] && !f[546];
	assign leaf[10355] = f[349] && !f[519] && f[436] && f[546];
	assign leaf[10356] = f[349] && f[519] && !f[375] && !f[295];
	assign leaf[10357] = f[349] && f[519] && !f[375] && f[295];
	assign leaf[10358] = f[349] && f[519] && f[375] && !f[579];
	assign leaf[10359] = f[349] && f[519] && f[375] && f[579];
	
	// Tree 749, Classifier 9, Iteration: 74
	assign leaf[10360] = !f[351] && !f[377] && !f[323] && !f[407];
	assign leaf[10361] = !f[351] && !f[377] && !f[323] && f[407];
	assign leaf[10362] = !f[351] && !f[377] && f[323] && !f[709];
	assign leaf[10363] = !f[351] && !f[377] && f[323] && f[709];
	assign leaf[10364] = !f[351] && f[377] && !f[652] && !f[713];
	assign leaf[10365] = !f[351] && f[377] && !f[652] && f[713];
	assign leaf[10366] = !f[351] && f[377] && f[652] && !f[412];
	assign leaf[10367] = !f[351] && f[377] && f[652] && f[412];
	assign leaf[10368] = f[351] && !f[511] && !f[434] && !f[152];
	assign leaf[10369] = f[351] && !f[511] && !f[434] && f[152];
	assign leaf[10370] = f[351] && !f[511] && f[434] && !f[320];
	assign leaf[10371] = f[351] && !f[511] && f[434] && f[320];
	assign leaf[10372] = f[351] && f[511] && !f[659] && !f[260];
	assign leaf[10373] = f[351] && f[511] && !f[659] && f[260];
	assign leaf[10374] = f[351] && f[511] && f[659] && !f[521];
	assign leaf[10375] = f[351] && f[511] && f[659] && f[521];
	
	// Tree 750, Classifier 0, Iteration: 75
	assign leaf[10376] = !f[602] && !f[576] && !f[460] && !f[205];
	assign leaf[10377] = !f[602] && !f[576] && !f[460] && f[205];
	assign leaf[10378] = !f[602] && !f[576] && f[460] && !f[351];
	assign leaf[10379] = !f[602] && !f[576] && f[460] && f[351];
	assign leaf[10380] = !f[602] && f[576] && !f[442] && !f[656];
	assign leaf[10381] = !f[602] && f[576] && !f[442] && f[656];
	assign leaf[10382] = !f[602] && f[576] && f[442];
	assign leaf[10383] = f[602] && !f[323] && !f[600] && !f[626];
	assign leaf[10384] = f[602] && !f[323] && !f[600] && f[626];
	assign leaf[10385] = f[602] && !f[323] && f[600] && !f[630];
	assign leaf[10386] = f[602] && !f[323] && f[600] && f[630];
	assign leaf[10387] = f[602] && f[323] && !f[264] && !f[433];
	assign leaf[10388] = f[602] && f[323] && !f[264] && f[433];
	assign leaf[10389] = f[602] && f[323] && f[264] && !f[626];
	assign leaf[10390] = f[602] && f[323] && f[264] && f[626];
	
	// Tree 751, Classifier 1, Iteration: 75
	assign leaf[10391] = !f[375] && !f[321] && !f[686] && !f[460];
	assign leaf[10392] = !f[375] && !f[321] && !f[686] && f[460];
	assign leaf[10393] = !f[375] && !f[321] && f[686] && !f[432];
	assign leaf[10394] = !f[375] && !f[321] && f[686] && f[432];
	assign leaf[10395] = !f[375] && f[321] && !f[213] && !f[269];
	assign leaf[10396] = !f[375] && f[321] && !f[213] && f[269];
	assign leaf[10397] = !f[375] && f[321] && f[213] && !f[460];
	assign leaf[10398] = !f[375] && f[321] && f[213] && f[460];
	assign leaf[10399] = f[375] && !f[321] && !f[403];
	assign leaf[10400] = f[375] && !f[321] && f[403];
	assign leaf[10401] = f[375] && f[321] && !f[687] && !f[129];
	assign leaf[10402] = f[375] && f[321] && !f[687] && f[129];
	assign leaf[10403] = f[375] && f[321] && f[687] && !f[377];
	assign leaf[10404] = f[375] && f[321] && f[687] && f[377];
	
	// Tree 752, Classifier 2, Iteration: 75
	assign leaf[10405] = !f[715] && !f[718] && !f[547] && !f[603];
	assign leaf[10406] = !f[715] && !f[718] && !f[547] && f[603];
	assign leaf[10407] = !f[715] && !f[718] && f[547] && !f[636];
	assign leaf[10408] = !f[715] && !f[718] && f[547] && f[636];
	assign leaf[10409] = !f[715] && f[718] && !f[492];
	assign leaf[10410] = !f[715] && f[718] && f[492];
	assign leaf[10411] = f[715] && !f[576] && !f[717];
	assign leaf[10412] = f[715] && !f[576] && f[717];
	assign leaf[10413] = f[715] && f[576] && !f[295];
	assign leaf[10414] = f[715] && f[576] && f[295];
	
	// Tree 753, Classifier 3, Iteration: 75
	assign leaf[10415] = !f[712] && !f[313] && !f[202] && !f[258];
	assign leaf[10416] = !f[712] && !f[313] && !f[202] && f[258];
	assign leaf[10417] = !f[712] && !f[313] && f[202] && !f[576];
	assign leaf[10418] = !f[712] && !f[313] && f[202] && f[576];
	assign leaf[10419] = !f[712] && f[313] && !f[525] && !f[685];
	assign leaf[10420] = !f[712] && f[313] && !f[525] && f[685];
	assign leaf[10421] = !f[712] && f[313] && f[525] && !f[397];
	assign leaf[10422] = !f[712] && f[313] && f[525] && f[397];
	assign leaf[10423] = f[712] && !f[684] && !f[178];
	assign leaf[10424] = f[712] && !f[684] && f[178];
	assign leaf[10425] = f[712] && f[684] && !f[576] && !f[356];
	assign leaf[10426] = f[712] && f[684] && !f[576] && f[356];
	assign leaf[10427] = f[712] && f[684] && f[576] && !f[299];
	assign leaf[10428] = f[712] && f[684] && f[576] && f[299];
	
	// Tree 754, Classifier 4, Iteration: 75
	assign leaf[10429] = !f[737] && !f[303] && !f[398] && !f[347];
	assign leaf[10430] = !f[737] && !f[303] && !f[398] && f[347];
	assign leaf[10431] = !f[737] && !f[303] && f[398] && !f[294];
	assign leaf[10432] = !f[737] && !f[303] && f[398] && f[294];
	assign leaf[10433] = !f[737] && f[303] && !f[453] && !f[324];
	assign leaf[10434] = !f[737] && f[303] && !f[453] && f[324];
	assign leaf[10435] = !f[737] && f[303] && f[453];
	assign leaf[10436] = f[737];
	
	// Tree 755, Classifier 5, Iteration: 75
	assign leaf[10437] = !f[402] && !f[484] && !f[631] && !f[493];
	assign leaf[10438] = !f[402] && !f[484] && !f[631] && f[493];
	assign leaf[10439] = !f[402] && !f[484] && f[631] && !f[601];
	assign leaf[10440] = !f[402] && !f[484] && f[631] && f[601];
	assign leaf[10441] = !f[402] && f[484] && !f[371] && !f[459];
	assign leaf[10442] = !f[402] && f[484] && !f[371] && f[459];
	assign leaf[10443] = !f[402] && f[484] && f[371] && !f[430];
	assign leaf[10444] = !f[402] && f[484] && f[371] && f[430];
	assign leaf[10445] = f[402] && !f[484] && !f[518] && !f[318];
	assign leaf[10446] = f[402] && !f[484] && !f[518] && f[318];
	assign leaf[10447] = f[402] && !f[484] && f[518] && !f[184];
	assign leaf[10448] = f[402] && !f[484] && f[518] && f[184];
	assign leaf[10449] = f[402] && f[484] && !f[625] && !f[317];
	assign leaf[10450] = f[402] && f[484] && !f[625] && f[317];
	assign leaf[10451] = f[402] && f[484] && f[625] && !f[489];
	assign leaf[10452] = f[402] && f[484] && f[625] && f[489];
	
	// Tree 756, Classifier 6, Iteration: 75
	assign leaf[10453] = !f[652] && !f[655] && !f[162] && !f[374];
	assign leaf[10454] = !f[652] && !f[655] && !f[162] && f[374];
	assign leaf[10455] = !f[652] && !f[655] && f[162] && !f[189];
	assign leaf[10456] = !f[652] && !f[655] && f[162] && f[189];
	assign leaf[10457] = !f[652] && f[655] && !f[241] && !f[211];
	assign leaf[10458] = !f[652] && f[655] && !f[241] && f[211];
	assign leaf[10459] = !f[652] && f[655] && f[241] && !f[379];
	assign leaf[10460] = !f[652] && f[655] && f[241] && f[379];
	assign leaf[10461] = f[652] && !f[488];
	assign leaf[10462] = f[652] && f[488];
	
	// Tree 757, Classifier 7, Iteration: 75
	assign leaf[10463] = !f[515] && !f[457] && !f[426] && !f[265];
	assign leaf[10464] = !f[515] && !f[457] && !f[426] && f[265];
	assign leaf[10465] = !f[515] && !f[457] && f[426] && !f[430];
	assign leaf[10466] = !f[515] && !f[457] && f[426] && f[430];
	assign leaf[10467] = !f[515] && f[457] && !f[460] && !f[569];
	assign leaf[10468] = !f[515] && f[457] && !f[460] && f[569];
	assign leaf[10469] = !f[515] && f[457] && f[460] && !f[372];
	assign leaf[10470] = !f[515] && f[457] && f[460] && f[372];
	assign leaf[10471] = f[515] && !f[428] && !f[426] && !f[291];
	assign leaf[10472] = f[515] && !f[428] && !f[426] && f[291];
	assign leaf[10473] = f[515] && !f[428] && f[426];
	assign leaf[10474] = f[515] && f[428] && !f[485] && !f[601];
	assign leaf[10475] = f[515] && f[428] && !f[485] && f[601];
	assign leaf[10476] = f[515] && f[428] && f[485] && !f[405];
	assign leaf[10477] = f[515] && f[428] && f[485] && f[405];
	
	// Tree 758, Classifier 8, Iteration: 75
	assign leaf[10478] = !f[186] && !f[129] && !f[151] && !f[266];
	assign leaf[10479] = !f[186] && !f[129] && !f[151] && f[266];
	assign leaf[10480] = !f[186] && !f[129] && f[151] && !f[576];
	assign leaf[10481] = !f[186] && !f[129] && f[151] && f[576];
	assign leaf[10482] = !f[186] && f[129] && !f[378] && !f[517];
	assign leaf[10483] = !f[186] && f[129] && !f[378] && f[517];
	assign leaf[10484] = !f[186] && f[129] && f[378] && !f[267];
	assign leaf[10485] = !f[186] && f[129] && f[378] && f[267];
	assign leaf[10486] = f[186] && !f[294] && !f[153] && !f[637];
	assign leaf[10487] = f[186] && !f[294] && !f[153] && f[637];
	assign leaf[10488] = f[186] && !f[294] && f[153] && !f[599];
	assign leaf[10489] = f[186] && !f[294] && f[153] && f[599];
	assign leaf[10490] = f[186] && f[294] && !f[348] && !f[319];
	assign leaf[10491] = f[186] && f[294] && !f[348] && f[319];
	assign leaf[10492] = f[186] && f[294] && f[348] && !f[262];
	assign leaf[10493] = f[186] && f[294] && f[348] && f[262];
	
	// Tree 759, Classifier 9, Iteration: 75
	assign leaf[10494] = !f[686] && !f[603] && !f[715] && !f[186];
	assign leaf[10495] = !f[686] && !f[603] && !f[715] && f[186];
	assign leaf[10496] = !f[686] && !f[603] && f[715] && !f[521];
	assign leaf[10497] = !f[686] && !f[603] && f[715] && f[521];
	assign leaf[10498] = !f[686] && f[603] && !f[181] && !f[744];
	assign leaf[10499] = !f[686] && f[603] && !f[181] && f[744];
	assign leaf[10500] = !f[686] && f[603] && f[181] && !f[659];
	assign leaf[10501] = !f[686] && f[603] && f[181] && f[659];
	assign leaf[10502] = f[686] && !f[572] && !f[518] && !f[547];
	assign leaf[10503] = f[686] && !f[572] && !f[518] && f[547];
	assign leaf[10504] = f[686] && !f[572] && f[518] && !f[264];
	assign leaf[10505] = f[686] && !f[572] && f[518] && f[264];
	assign leaf[10506] = f[686] && f[572] && !f[428] && !f[489];
	assign leaf[10507] = f[686] && f[572] && !f[428] && f[489];
	assign leaf[10508] = f[686] && f[572] && f[428] && !f[604];
	assign leaf[10509] = f[686] && f[572] && f[428] && f[604];
	
	// Tree 760, Classifier 0, Iteration: 76
	assign leaf[10510] = !f[213] && !f[544] && !f[384] && !f[408];
	assign leaf[10511] = !f[213] && !f[544] && !f[384] && f[408];
	assign leaf[10512] = !f[213] && !f[544] && f[384] && !f[215];
	assign leaf[10513] = !f[213] && !f[544] && f[384] && f[215];
	assign leaf[10514] = !f[213] && f[544] && !f[296] && !f[481];
	assign leaf[10515] = !f[213] && f[544] && !f[296] && f[481];
	assign leaf[10516] = !f[213] && f[544] && f[296] && !f[494];
	assign leaf[10517] = !f[213] && f[544] && f[296] && f[494];
	assign leaf[10518] = f[213] && !f[323] && !f[347] && !f[519];
	assign leaf[10519] = f[213] && !f[323] && !f[347] && f[519];
	assign leaf[10520] = f[213] && !f[323] && f[347] && !f[316];
	assign leaf[10521] = f[213] && !f[323] && f[347] && f[316];
	assign leaf[10522] = f[213] && f[323] && !f[153] && !f[428];
	assign leaf[10523] = f[213] && f[323] && !f[153] && f[428];
	assign leaf[10524] = f[213] && f[323] && f[153] && !f[490];
	assign leaf[10525] = f[213] && f[323] && f[153] && f[490];
	
	// Tree 761, Classifier 1, Iteration: 76
	assign leaf[10526] = !f[715] && !f[401] && !f[376] && !f[153];
	assign leaf[10527] = !f[715] && !f[401] && !f[376] && f[153];
	assign leaf[10528] = !f[715] && !f[401] && f[376] && !f[658];
	assign leaf[10529] = !f[715] && !f[401] && f[376] && f[658];
	assign leaf[10530] = !f[715] && f[401] && !f[461] && !f[345];
	assign leaf[10531] = !f[715] && f[401] && !f[461] && f[345];
	assign leaf[10532] = !f[715] && f[401] && f[461];
	assign leaf[10533] = f[715] && !f[403];
	assign leaf[10534] = f[715] && f[403];
	
	// Tree 762, Classifier 2, Iteration: 76
	assign leaf[10535] = !f[258] && !f[636] && !f[553] && !f[470];
	assign leaf[10536] = !f[258] && !f[636] && !f[553] && f[470];
	assign leaf[10537] = !f[258] && !f[636] && f[553] && !f[607];
	assign leaf[10538] = !f[258] && !f[636] && f[553] && f[607];
	assign leaf[10539] = !f[258] && f[636] && !f[524] && !f[260];
	assign leaf[10540] = !f[258] && f[636] && !f[524] && f[260];
	assign leaf[10541] = !f[258] && f[636] && f[524] && !f[577];
	assign leaf[10542] = !f[258] && f[636] && f[524] && f[577];
	assign leaf[10543] = f[258] && !f[455] && !f[635] && !f[244];
	assign leaf[10544] = f[258] && !f[455] && !f[635] && f[244];
	assign leaf[10545] = f[258] && !f[455] && f[635] && !f[604];
	assign leaf[10546] = f[258] && !f[455] && f[635] && f[604];
	assign leaf[10547] = f[258] && f[455];
	
	// Tree 763, Classifier 3, Iteration: 76
	assign leaf[10548] = !f[708] && !f[466] && !f[718] && !f[200];
	assign leaf[10549] = !f[708] && !f[466] && !f[718] && f[200];
	assign leaf[10550] = !f[708] && !f[466] && f[718] && !f[213];
	assign leaf[10551] = !f[708] && !f[466] && f[718] && f[213];
	assign leaf[10552] = !f[708] && f[466] && !f[355] && !f[403];
	assign leaf[10553] = !f[708] && f[466] && !f[355] && f[403];
	assign leaf[10554] = !f[708] && f[466] && f[355] && !f[543];
	assign leaf[10555] = !f[708] && f[466] && f[355] && f[543];
	assign leaf[10556] = f[708] && !f[599] && !f[491];
	assign leaf[10557] = f[708] && !f[599] && f[491];
	assign leaf[10558] = f[708] && f[599];
	
	// Tree 764, Classifier 4, Iteration: 76
	assign leaf[10559] = !f[746] && !f[376] && !f[321] && !f[182];
	assign leaf[10560] = !f[746] && !f[376] && !f[321] && f[182];
	assign leaf[10561] = !f[746] && !f[376] && f[321] && !f[238];
	assign leaf[10562] = !f[746] && !f[376] && f[321] && f[238];
	assign leaf[10563] = !f[746] && f[376] && !f[435] && !f[296];
	assign leaf[10564] = !f[746] && f[376] && !f[435] && f[296];
	assign leaf[10565] = !f[746] && f[376] && f[435] && !f[155];
	assign leaf[10566] = !f[746] && f[376] && f[435] && f[155];
	assign leaf[10567] = f[746];
	
	// Tree 765, Classifier 5, Iteration: 76
	assign leaf[10568] = !f[707] && !f[402] && !f[243] && !f[187];
	assign leaf[10569] = !f[707] && !f[402] && !f[243] && f[187];
	assign leaf[10570] = !f[707] && !f[402] && f[243] && !f[240];
	assign leaf[10571] = !f[707] && !f[402] && f[243] && f[240];
	assign leaf[10572] = !f[707] && f[402] && !f[156] && !f[177];
	assign leaf[10573] = !f[707] && f[402] && !f[156] && f[177];
	assign leaf[10574] = !f[707] && f[402] && f[156] && !f[270];
	assign leaf[10575] = !f[707] && f[402] && f[156] && f[270];
	assign leaf[10576] = f[707] && !f[627];
	assign leaf[10577] = f[707] && f[627];
	
	// Tree 766, Classifier 6, Iteration: 76
	assign leaf[10578] = !f[682] && !f[638] && !f[610] && !f[406];
	assign leaf[10579] = !f[682] && !f[638] && !f[610] && f[406];
	assign leaf[10580] = !f[682] && !f[638] && f[610] && !f[315];
	assign leaf[10581] = !f[682] && !f[638] && f[610] && f[315];
	assign leaf[10582] = !f[682] && f[638];
	assign leaf[10583] = f[682];
	
	// Tree 767, Classifier 7, Iteration: 76
	assign leaf[10584] = !f[510] && !f[464] && !f[547] && !f[176];
	assign leaf[10585] = !f[510] && !f[464] && !f[547] && f[176];
	assign leaf[10586] = !f[510] && !f[464] && f[547] && !f[377];
	assign leaf[10587] = !f[510] && !f[464] && f[547] && f[377];
	assign leaf[10588] = !f[510] && f[464] && !f[383] && !f[518];
	assign leaf[10589] = !f[510] && f[464] && !f[383] && f[518];
	assign leaf[10590] = !f[510] && f[464] && f[383] && !f[326];
	assign leaf[10591] = !f[510] && f[464] && f[383] && f[326];
	assign leaf[10592] = f[510] && !f[685] && !f[661] && !f[314];
	assign leaf[10593] = f[510] && !f[685] && !f[661] && f[314];
	assign leaf[10594] = f[510] && !f[685] && f[661];
	assign leaf[10595] = f[510] && f[685] && !f[296];
	assign leaf[10596] = f[510] && f[685] && f[296];
	
	// Tree 768, Classifier 8, Iteration: 76
	assign leaf[10597] = !f[236] && !f[260] && !f[262] && !f[238];
	assign leaf[10598] = !f[236] && !f[260] && !f[262] && f[238];
	assign leaf[10599] = !f[236] && !f[260] && f[262] && !f[240];
	assign leaf[10600] = !f[236] && !f[260] && f[262] && f[240];
	assign leaf[10601] = !f[236] && f[260] && !f[316] && !f[596];
	assign leaf[10602] = !f[236] && f[260] && !f[316] && f[596];
	assign leaf[10603] = !f[236] && f[260] && f[316] && !f[271];
	assign leaf[10604] = !f[236] && f[260] && f[316] && f[271];
	assign leaf[10605] = f[236] && !f[204] && !f[319] && !f[293];
	assign leaf[10606] = f[236] && !f[204] && !f[319] && f[293];
	assign leaf[10607] = f[236] && !f[204] && f[319] && !f[293];
	assign leaf[10608] = f[236] && !f[204] && f[319] && f[293];
	assign leaf[10609] = f[236] && f[204] && !f[352] && !f[488];
	assign leaf[10610] = f[236] && f[204] && !f[352] && f[488];
	assign leaf[10611] = f[236] && f[204] && f[352] && !f[300];
	assign leaf[10612] = f[236] && f[204] && f[352] && f[300];
	
	// Tree 769, Classifier 9, Iteration: 76
	assign leaf[10613] = !f[742] && !f[162] && !f[229] && !f[740];
	assign leaf[10614] = !f[742] && !f[162] && !f[229] && f[740];
	assign leaf[10615] = !f[742] && !f[162] && f[229] && !f[260];
	assign leaf[10616] = !f[742] && !f[162] && f[229] && f[260];
	assign leaf[10617] = !f[742] && f[162] && !f[246];
	assign leaf[10618] = !f[742] && f[162] && f[246];
	assign leaf[10619] = f[742] && !f[328] && !f[259] && !f[326];
	assign leaf[10620] = f[742] && !f[328] && !f[259] && f[326];
	assign leaf[10621] = f[742] && !f[328] && f[259];
	assign leaf[10622] = f[742] && f[328] && !f[345];
	assign leaf[10623] = f[742] && f[328] && f[345] && !f[494];
	assign leaf[10624] = f[742] && f[328] && f[345] && f[494];
	
	// Tree 770, Classifier 0, Iteration: 77
	assign leaf[10625] = !f[434] && !f[486] && !f[489] && !f[276];
	assign leaf[10626] = !f[434] && !f[486] && !f[489] && f[276];
	assign leaf[10627] = !f[434] && !f[486] && f[489] && !f[354];
	assign leaf[10628] = !f[434] && !f[486] && f[489] && f[354];
	assign leaf[10629] = !f[434] && f[486] && !f[287] && !f[489];
	assign leaf[10630] = !f[434] && f[486] && !f[287] && f[489];
	assign leaf[10631] = !f[434] && f[486] && f[287] && !f[291];
	assign leaf[10632] = !f[434] && f[486] && f[287] && f[291];
	assign leaf[10633] = f[434] && !f[357] && !f[461];
	assign leaf[10634] = f[434] && !f[357] && f[461];
	assign leaf[10635] = f[434] && f[357] && !f[158] && !f[546];
	assign leaf[10636] = f[434] && f[357] && !f[158] && f[546];
	assign leaf[10637] = f[434] && f[357] && f[158] && !f[409];
	assign leaf[10638] = f[434] && f[357] && f[158] && f[409];
	
	// Tree 771, Classifier 1, Iteration: 77
	assign leaf[10639] = !f[384] && !f[131] && !f[270] && !f[187];
	assign leaf[10640] = !f[384] && !f[131] && !f[270] && f[187];
	assign leaf[10641] = !f[384] && !f[131] && f[270] && !f[408];
	assign leaf[10642] = !f[384] && !f[131] && f[270] && f[408];
	assign leaf[10643] = !f[384] && f[131] && !f[324] && !f[129];
	assign leaf[10644] = !f[384] && f[131] && !f[324] && f[129];
	assign leaf[10645] = !f[384] && f[131] && f[324] && !f[241];
	assign leaf[10646] = !f[384] && f[131] && f[324] && f[241];
	assign leaf[10647] = f[384];
	
	// Tree 772, Classifier 2, Iteration: 77
	assign leaf[10648] = !f[125] && !f[546] && !f[657] && !f[688];
	assign leaf[10649] = !f[125] && !f[546] && !f[657] && f[688];
	assign leaf[10650] = !f[125] && !f[546] && f[657] && !f[376];
	assign leaf[10651] = !f[125] && !f[546] && f[657] && f[376];
	assign leaf[10652] = !f[125] && f[546] && !f[219] && !f[711];
	assign leaf[10653] = !f[125] && f[546] && !f[219] && f[711];
	assign leaf[10654] = !f[125] && f[546] && f[219] && !f[564];
	assign leaf[10655] = !f[125] && f[546] && f[219] && f[564];
	assign leaf[10656] = f[125] && !f[240] && !f[381] && !f[300];
	assign leaf[10657] = f[125] && !f[240] && !f[381] && f[300];
	assign leaf[10658] = f[125] && !f[240] && f[381] && !f[243];
	assign leaf[10659] = f[125] && !f[240] && f[381] && f[243];
	assign leaf[10660] = f[125] && f[240] && !f[438] && !f[499];
	assign leaf[10661] = f[125] && f[240] && !f[438] && f[499];
	assign leaf[10662] = f[125] && f[240] && f[438] && !f[266];
	assign leaf[10663] = f[125] && f[240] && f[438] && f[266];
	
	// Tree 773, Classifier 3, Iteration: 77
	assign leaf[10664] = !f[427] && !f[651] && !f[712] && !f[626];
	assign leaf[10665] = !f[427] && !f[651] && !f[712] && f[626];
	assign leaf[10666] = !f[427] && !f[651] && f[712] && !f[488];
	assign leaf[10667] = !f[427] && !f[651] && f[712] && f[488];
	assign leaf[10668] = !f[427] && f[651] && !f[542] && !f[461];
	assign leaf[10669] = !f[427] && f[651] && !f[542] && f[461];
	assign leaf[10670] = !f[427] && f[651] && f[542] && !f[656];
	assign leaf[10671] = !f[427] && f[651] && f[542] && f[656];
	assign leaf[10672] = f[427] && !f[436] && !f[236] && !f[295];
	assign leaf[10673] = f[427] && !f[436] && !f[236] && f[295];
	assign leaf[10674] = f[427] && !f[436] && f[236] && !f[597];
	assign leaf[10675] = f[427] && !f[436] && f[236] && f[597];
	assign leaf[10676] = f[427] && f[436] && !f[580] && !f[568];
	assign leaf[10677] = f[427] && f[436] && !f[580] && f[568];
	assign leaf[10678] = f[427] && f[436] && f[580] && !f[658];
	assign leaf[10679] = f[427] && f[436] && f[580] && f[658];
	
	// Tree 774, Classifier 4, Iteration: 77
	assign leaf[10680] = !f[465] && !f[238] && !f[213] && !f[215];
	assign leaf[10681] = !f[465] && !f[238] && !f[213] && f[215];
	assign leaf[10682] = !f[465] && !f[238] && f[213] && !f[182];
	assign leaf[10683] = !f[465] && !f[238] && f[213] && f[182];
	assign leaf[10684] = !f[465] && f[238] && !f[240] && !f[186];
	assign leaf[10685] = !f[465] && f[238] && !f[240] && f[186];
	assign leaf[10686] = !f[465] && f[238] && f[240] && !f[242];
	assign leaf[10687] = !f[465] && f[238] && f[240] && f[242];
	assign leaf[10688] = f[465] && !f[340] && !f[242] && !f[328];
	assign leaf[10689] = f[465] && !f[340] && !f[242] && f[328];
	assign leaf[10690] = f[465] && !f[340] && f[242] && !f[328];
	assign leaf[10691] = f[465] && !f[340] && f[242] && f[328];
	assign leaf[10692] = f[465] && f[340] && !f[240] && !f[352];
	assign leaf[10693] = f[465] && f[340] && !f[240] && f[352];
	assign leaf[10694] = f[465] && f[340] && f[240];
	
	// Tree 775, Classifier 5, Iteration: 77
	assign leaf[10695] = !f[190] && !f[130] && !f[406] && !f[464];
	assign leaf[10696] = !f[190] && !f[130] && !f[406] && f[464];
	assign leaf[10697] = !f[190] && !f[130] && f[406] && !f[325];
	assign leaf[10698] = !f[190] && !f[130] && f[406] && f[325];
	assign leaf[10699] = !f[190] && f[130] && !f[215] && !f[154];
	assign leaf[10700] = !f[190] && f[130] && !f[215] && f[154];
	assign leaf[10701] = !f[190] && f[130] && f[215] && !f[239];
	assign leaf[10702] = !f[190] && f[130] && f[215] && f[239];
	assign leaf[10703] = f[190] && !f[214] && !f[540] && !f[492];
	assign leaf[10704] = f[190] && !f[214] && !f[540] && f[492];
	assign leaf[10705] = f[190] && !f[214] && f[540] && !f[625];
	assign leaf[10706] = f[190] && !f[214] && f[540] && f[625];
	assign leaf[10707] = f[190] && f[214] && !f[275] && !f[160];
	assign leaf[10708] = f[190] && f[214] && !f[275] && f[160];
	assign leaf[10709] = f[190] && f[214] && f[275] && !f[270];
	assign leaf[10710] = f[190] && f[214] && f[275] && f[270];
	
	// Tree 776, Classifier 6, Iteration: 77
	assign leaf[10711] = !f[214] && !f[637] && !f[295] && !f[247];
	assign leaf[10712] = !f[214] && !f[637] && !f[295] && f[247];
	assign leaf[10713] = !f[214] && !f[637] && f[295] && !f[265];
	assign leaf[10714] = !f[214] && !f[637] && f[295] && f[265];
	assign leaf[10715] = !f[214] && f[637];
	assign leaf[10716] = f[214] && !f[348] && !f[377] && !f[320];
	assign leaf[10717] = f[214] && !f[348] && !f[377] && f[320];
	assign leaf[10718] = f[214] && !f[348] && f[377] && !f[316];
	assign leaf[10719] = f[214] && !f[348] && f[377] && f[316];
	assign leaf[10720] = f[214] && f[348] && !f[687] && !f[235];
	assign leaf[10721] = f[214] && f[348] && !f[687] && f[235];
	assign leaf[10722] = f[214] && f[348] && f[687];
	
	// Tree 777, Classifier 7, Iteration: 77
	assign leaf[10723] = !f[528] && !f[527] && !f[709] && !f[708];
	assign leaf[10724] = !f[528] && !f[527] && !f[709] && f[708];
	assign leaf[10725] = !f[528] && !f[527] && f[709] && !f[630];
	assign leaf[10726] = !f[528] && !f[527] && f[709] && f[630];
	assign leaf[10727] = !f[528] && f[527] && !f[242];
	assign leaf[10728] = !f[528] && f[527] && f[242];
	assign leaf[10729] = f[528] && !f[600];
	assign leaf[10730] = f[528] && f[600];
	
	// Tree 778, Classifier 8, Iteration: 77
	assign leaf[10731] = !f[135] && !f[328] && !f[405] && !f[430];
	assign leaf[10732] = !f[135] && !f[328] && !f[405] && f[430];
	assign leaf[10733] = !f[135] && !f[328] && f[405] && !f[656];
	assign leaf[10734] = !f[135] && !f[328] && f[405] && f[656];
	assign leaf[10735] = !f[135] && f[328] && !f[458] && !f[298];
	assign leaf[10736] = !f[135] && f[328] && !f[458] && f[298];
	assign leaf[10737] = !f[135] && f[328] && f[458] && !f[405];
	assign leaf[10738] = !f[135] && f[328] && f[458] && f[405];
	assign leaf[10739] = f[135] && !f[270];
	assign leaf[10740] = f[135] && f[270];
	
	// Tree 779, Classifier 9, Iteration: 77
	assign leaf[10741] = !f[350] && !f[384] && !f[467] && !f[378];
	assign leaf[10742] = !f[350] && !f[384] && !f[467] && f[378];
	assign leaf[10743] = !f[350] && !f[384] && f[467] && !f[288];
	assign leaf[10744] = !f[350] && !f[384] && f[467] && f[288];
	assign leaf[10745] = !f[350] && f[384] && !f[467] && !f[215];
	assign leaf[10746] = !f[350] && f[384] && !f[467] && f[215];
	assign leaf[10747] = !f[350] && f[384] && f[467] && !f[246];
	assign leaf[10748] = !f[350] && f[384] && f[467] && f[246];
	assign leaf[10749] = f[350] && !f[324] && !f[651] && !f[352];
	assign leaf[10750] = f[350] && !f[324] && !f[651] && f[352];
	assign leaf[10751] = f[350] && !f[324] && f[651];
	assign leaf[10752] = f[350] && f[324] && !f[487] && !f[384];
	assign leaf[10753] = f[350] && f[324] && !f[487] && f[384];
	assign leaf[10754] = f[350] && f[324] && f[487] && !f[628];
	assign leaf[10755] = f[350] && f[324] && f[487] && f[628];
	
	// Tree 780, Classifier 0, Iteration: 78
	assign leaf[10756] = !f[512] && !f[462] && !f[597] && !f[155];
	assign leaf[10757] = !f[512] && !f[462] && !f[597] && f[155];
	assign leaf[10758] = !f[512] && !f[462] && f[597] && !f[606];
	assign leaf[10759] = !f[512] && !f[462] && f[597] && f[606];
	assign leaf[10760] = !f[512] && f[462] && !f[481];
	assign leaf[10761] = !f[512] && f[462] && f[481];
	assign leaf[10762] = f[512] && !f[654] && !f[575] && !f[484];
	assign leaf[10763] = f[512] && !f[654] && !f[575] && f[484];
	assign leaf[10764] = f[512] && !f[654] && f[575] && !f[437];
	assign leaf[10765] = f[512] && !f[654] && f[575] && f[437];
	assign leaf[10766] = f[512] && f[654] && !f[247] && !f[400];
	assign leaf[10767] = f[512] && f[654] && !f[247] && f[400];
	assign leaf[10768] = f[512] && f[654] && f[247];
	
	// Tree 781, Classifier 1, Iteration: 78
	assign leaf[10769] = !f[316] && !f[635] && !f[566] && !f[540];
	assign leaf[10770] = !f[316] && !f[635] && !f[566] && f[540];
	assign leaf[10771] = !f[316] && !f[635] && f[566] && !f[404];
	assign leaf[10772] = !f[316] && !f[635] && f[566] && f[404];
	assign leaf[10773] = !f[316] && f[635] && !f[516] && !f[267];
	assign leaf[10774] = !f[316] && f[635] && !f[516] && f[267];
	assign leaf[10775] = !f[316] && f[635] && f[516] && !f[152];
	assign leaf[10776] = !f[316] && f[635] && f[516] && f[152];
	assign leaf[10777] = f[316] && !f[598];
	assign leaf[10778] = f[316] && f[598];
	
	// Tree 782, Classifier 2, Iteration: 78
	assign leaf[10779] = !f[501] && !f[570] && !f[539] && !f[356];
	assign leaf[10780] = !f[501] && !f[570] && !f[539] && f[356];
	assign leaf[10781] = !f[501] && !f[570] && f[539] && !f[459];
	assign leaf[10782] = !f[501] && !f[570] && f[539] && f[459];
	assign leaf[10783] = !f[501] && f[570] && !f[406] && !f[524];
	assign leaf[10784] = !f[501] && f[570] && !f[406] && f[524];
	assign leaf[10785] = !f[501] && f[570] && f[406] && !f[273];
	assign leaf[10786] = !f[501] && f[570] && f[406] && f[273];
	assign leaf[10787] = f[501] && !f[322];
	assign leaf[10788] = f[501] && f[322];
	
	// Tree 783, Classifier 3, Iteration: 78
	assign leaf[10789] = !f[384] && !f[487] && !f[124] && !f[554];
	assign leaf[10790] = !f[384] && !f[487] && !f[124] && f[554];
	assign leaf[10791] = !f[384] && !f[487] && f[124] && !f[207];
	assign leaf[10792] = !f[384] && !f[487] && f[124] && f[207];
	assign leaf[10793] = !f[384] && f[487] && !f[570] && !f[294];
	assign leaf[10794] = !f[384] && f[487] && !f[570] && f[294];
	assign leaf[10795] = !f[384] && f[487] && f[570] && !f[460];
	assign leaf[10796] = !f[384] && f[487] && f[570] && f[460];
	assign leaf[10797] = f[384] && !f[295] && !f[439] && !f[496];
	assign leaf[10798] = f[384] && !f[295] && !f[439] && f[496];
	assign leaf[10799] = f[384] && !f[295] && f[439] && !f[158];
	assign leaf[10800] = f[384] && !f[295] && f[439] && f[158];
	assign leaf[10801] = f[384] && f[295] && !f[239] && !f[261];
	assign leaf[10802] = f[384] && f[295] && !f[239] && f[261];
	assign leaf[10803] = f[384] && f[295] && f[239] && !f[126];
	assign leaf[10804] = f[384] && f[295] && f[239] && f[126];
	
	// Tree 784, Classifier 4, Iteration: 78
	assign leaf[10805] = !f[102] && !f[430] && !f[379] && !f[580];
	assign leaf[10806] = !f[102] && !f[430] && !f[379] && f[580];
	assign leaf[10807] = !f[102] && !f[430] && f[379] && !f[459];
	assign leaf[10808] = !f[102] && !f[430] && f[379] && f[459];
	assign leaf[10809] = !f[102] && f[430] && !f[709] && !f[579];
	assign leaf[10810] = !f[102] && f[430] && !f[709] && f[579];
	assign leaf[10811] = !f[102] && f[430] && f[709] && !f[570];
	assign leaf[10812] = !f[102] && f[430] && f[709] && f[570];
	assign leaf[10813] = f[102] && !f[185];
	assign leaf[10814] = f[102] && f[185];
	
	// Tree 785, Classifier 5, Iteration: 78
	assign leaf[10815] = !f[99] && !f[153] && !f[102] && !f[687];
	assign leaf[10816] = !f[99] && !f[153] && !f[102] && f[687];
	assign leaf[10817] = !f[99] && !f[153] && f[102] && !f[464];
	assign leaf[10818] = !f[99] && !f[153] && f[102] && f[464];
	assign leaf[10819] = !f[99] && f[153] && !f[263] && !f[268];
	assign leaf[10820] = !f[99] && f[153] && !f[263] && f[268];
	assign leaf[10821] = !f[99] && f[153] && f[263] && !f[373];
	assign leaf[10822] = !f[99] && f[153] && f[263] && f[373];
	assign leaf[10823] = f[99] && !f[181] && !f[294] && !f[289];
	assign leaf[10824] = f[99] && !f[181] && !f[294] && f[289];
	assign leaf[10825] = f[99] && !f[181] && f[294];
	assign leaf[10826] = f[99] && f[181] && !f[458] && !f[237];
	assign leaf[10827] = f[99] && f[181] && !f[458] && f[237];
	assign leaf[10828] = f[99] && f[181] && f[458];
	
	// Tree 786, Classifier 6, Iteration: 78
	assign leaf[10829] = !f[571] && !f[574] && !f[541] && !f[578];
	assign leaf[10830] = !f[571] && !f[574] && !f[541] && f[578];
	assign leaf[10831] = !f[571] && !f[574] && f[541] && !f[384];
	assign leaf[10832] = !f[571] && !f[574] && f[541] && f[384];
	assign leaf[10833] = !f[571] && f[574] && !f[156] && !f[270];
	assign leaf[10834] = !f[571] && f[574] && !f[156] && f[270];
	assign leaf[10835] = !f[571] && f[574] && f[156] && !f[100];
	assign leaf[10836] = !f[571] && f[574] && f[156] && f[100];
	assign leaf[10837] = f[571] && !f[486] && !f[426] && !f[262];
	assign leaf[10838] = f[571] && !f[486] && !f[426] && f[262];
	assign leaf[10839] = f[571] && !f[486] && f[426] && !f[272];
	assign leaf[10840] = f[571] && !f[486] && f[426] && f[272];
	assign leaf[10841] = f[571] && f[486] && !f[540] && !f[514];
	assign leaf[10842] = f[571] && f[486] && !f[540] && f[514];
	assign leaf[10843] = f[571] && f[486] && f[540] && !f[400];
	assign leaf[10844] = f[571] && f[486] && f[540] && f[400];
	
	// Tree 787, Classifier 7, Iteration: 78
	assign leaf[10845] = !f[452] && !f[577] && !f[689] && !f[180];
	assign leaf[10846] = !f[452] && !f[577] && !f[689] && f[180];
	assign leaf[10847] = !f[452] && !f[577] && f[689] && !f[686];
	assign leaf[10848] = !f[452] && !f[577] && f[689] && f[686];
	assign leaf[10849] = !f[452] && f[577] && !f[626] && !f[202];
	assign leaf[10850] = !f[452] && f[577] && !f[626] && f[202];
	assign leaf[10851] = !f[452] && f[577] && f[626] && !f[157];
	assign leaf[10852] = !f[452] && f[577] && f[626] && f[157];
	assign leaf[10853] = f[452] && !f[427];
	assign leaf[10854] = f[452] && f[427];
	
	// Tree 788, Classifier 8, Iteration: 78
	assign leaf[10855] = !f[508] && !f[399] && !f[276] && !f[549];
	assign leaf[10856] = !f[508] && !f[399] && !f[276] && f[549];
	assign leaf[10857] = !f[508] && !f[399] && f[276] && !f[298];
	assign leaf[10858] = !f[508] && !f[399] && f[276] && f[298];
	assign leaf[10859] = !f[508] && f[399] && !f[346] && !f[353];
	assign leaf[10860] = !f[508] && f[399] && !f[346] && f[353];
	assign leaf[10861] = !f[508] && f[399] && f[346] && !f[432];
	assign leaf[10862] = !f[508] && f[399] && f[346] && f[432];
	assign leaf[10863] = f[508] && !f[538];
	assign leaf[10864] = f[508] && f[538];
	
	// Tree 789, Classifier 9, Iteration: 78
	assign leaf[10865] = !f[575] && !f[294] && !f[685] && !f[345];
	assign leaf[10866] = !f[575] && !f[294] && !f[685] && f[345];
	assign leaf[10867] = !f[575] && !f[294] && f[685] && !f[520];
	assign leaf[10868] = !f[575] && !f[294] && f[685] && f[520];
	assign leaf[10869] = !f[575] && f[294] && !f[301] && !f[259];
	assign leaf[10870] = !f[575] && f[294] && !f[301] && f[259];
	assign leaf[10871] = !f[575] && f[294] && f[301] && !f[433];
	assign leaf[10872] = !f[575] && f[294] && f[301] && f[433];
	assign leaf[10873] = f[575] && !f[517] && !f[209] && !f[181];
	assign leaf[10874] = f[575] && !f[517] && !f[209] && f[181];
	assign leaf[10875] = f[575] && !f[517] && f[209] && !f[456];
	assign leaf[10876] = f[575] && !f[517] && f[209] && f[456];
	assign leaf[10877] = f[575] && f[517] && !f[456] && !f[458];
	assign leaf[10878] = f[575] && f[517] && !f[456] && f[458];
	assign leaf[10879] = f[575] && f[517] && f[456] && !f[657];
	assign leaf[10880] = f[575] && f[517] && f[456] && f[657];
	
	// Tree 790, Classifier 0, Iteration: 79
	assign leaf[10881] = !f[607] && !f[688] && !f[192] && !f[258];
	assign leaf[10882] = !f[607] && !f[688] && !f[192] && f[258];
	assign leaf[10883] = !f[607] && !f[688] && f[192];
	assign leaf[10884] = !f[607] && f[688];
	assign leaf[10885] = f[607] && !f[633] && !f[439];
	assign leaf[10886] = f[607] && !f[633] && f[439];
	assign leaf[10887] = f[607] && f[633] && !f[208] && !f[371];
	assign leaf[10888] = f[607] && f[633] && !f[208] && f[371];
	assign leaf[10889] = f[607] && f[633] && f[208] && !f[157];
	assign leaf[10890] = f[607] && f[633] && f[208] && f[157];
	
	// Tree 791, Classifier 1, Iteration: 79
	assign leaf[10891] = !f[603] && !f[209] && !f[265] && !f[346];
	assign leaf[10892] = !f[603] && !f[209] && !f[265] && f[346];
	assign leaf[10893] = !f[603] && !f[209] && f[265] && !f[636];
	assign leaf[10894] = !f[603] && !f[209] && f[265] && f[636];
	assign leaf[10895] = !f[603] && f[209] && !f[238] && !f[295];
	assign leaf[10896] = !f[603] && f[209] && !f[238] && f[295];
	assign leaf[10897] = !f[603] && f[209] && f[238] && !f[325];
	assign leaf[10898] = !f[603] && f[209] && f[238] && f[325];
	assign leaf[10899] = f[603] && !f[546] && !f[578] && !f[210];
	assign leaf[10900] = f[603] && !f[546] && !f[578] && f[210];
	assign leaf[10901] = f[603] && !f[546] && f[578] && !f[492];
	assign leaf[10902] = f[603] && !f[546] && f[578] && f[492];
	assign leaf[10903] = f[603] && f[546] && !f[241] && !f[158];
	assign leaf[10904] = f[603] && f[546] && !f[241] && f[158];
	assign leaf[10905] = f[603] && f[546] && f[241] && !f[129];
	assign leaf[10906] = f[603] && f[546] && f[241] && f[129];
	
	// Tree 792, Classifier 2, Iteration: 79
	assign leaf[10907] = !f[622] && !f[216] && !f[102] && !f[633];
	assign leaf[10908] = !f[622] && !f[216] && !f[102] && f[633];
	assign leaf[10909] = !f[622] && !f[216] && f[102] && !f[601];
	assign leaf[10910] = !f[622] && !f[216] && f[102] && f[601];
	assign leaf[10911] = !f[622] && f[216] && !f[600] && !f[536];
	assign leaf[10912] = !f[622] && f[216] && !f[600] && f[536];
	assign leaf[10913] = !f[622] && f[216] && f[600] && !f[662];
	assign leaf[10914] = !f[622] && f[216] && f[600] && f[662];
	assign leaf[10915] = f[622] && !f[634] && !f[551] && !f[352];
	assign leaf[10916] = f[622] && !f[634] && !f[551] && f[352];
	assign leaf[10917] = f[622] && !f[634] && f[551] && !f[544];
	assign leaf[10918] = f[622] && !f[634] && f[551] && f[544];
	assign leaf[10919] = f[622] && f[634] && !f[271];
	assign leaf[10920] = f[622] && f[634] && f[271];
	
	// Tree 793, Classifier 3, Iteration: 79
	assign leaf[10921] = !f[346] && !f[433] && !f[462] && !f[314];
	assign leaf[10922] = !f[346] && !f[433] && !f[462] && f[314];
	assign leaf[10923] = !f[346] && !f[433] && f[462] && !f[298];
	assign leaf[10924] = !f[346] && !f[433] && f[462] && f[298];
	assign leaf[10925] = !f[346] && f[433] && !f[321] && !f[372];
	assign leaf[10926] = !f[346] && f[433] && !f[321] && f[372];
	assign leaf[10927] = !f[346] && f[433] && f[321] && !f[180];
	assign leaf[10928] = !f[346] && f[433] && f[321] && f[180];
	assign leaf[10929] = f[346] && !f[470] && !f[375] && !f[378];
	assign leaf[10930] = f[346] && !f[470] && !f[375] && f[378];
	assign leaf[10931] = f[346] && !f[470] && f[375] && !f[289];
	assign leaf[10932] = f[346] && !f[470] && f[375] && f[289];
	assign leaf[10933] = f[346] && f[470] && !f[463] && !f[410];
	assign leaf[10934] = f[346] && f[470] && !f[463] && f[410];
	assign leaf[10935] = f[346] && f[470] && f[463];
	
	// Tree 794, Classifier 4, Iteration: 79
	assign leaf[10936] = !f[685] && !f[320] && !f[289] && !f[287];
	assign leaf[10937] = !f[685] && !f[320] && !f[289] && f[287];
	assign leaf[10938] = !f[685] && !f[320] && f[289] && !f[180];
	assign leaf[10939] = !f[685] && !f[320] && f[289] && f[180];
	assign leaf[10940] = !f[685] && f[320] && !f[237] && !f[211];
	assign leaf[10941] = !f[685] && f[320] && !f[237] && f[211];
	assign leaf[10942] = !f[685] && f[320] && f[237] && !f[289];
	assign leaf[10943] = !f[685] && f[320] && f[237] && f[289];
	assign leaf[10944] = f[685] && !f[239] && !f[184] && !f[322];
	assign leaf[10945] = f[685] && !f[239] && !f[184] && f[322];
	assign leaf[10946] = f[685] && !f[239] && f[184] && !f[183];
	assign leaf[10947] = f[685] && !f[239] && f[184] && f[183];
	assign leaf[10948] = f[685] && f[239] && !f[322] && !f[433];
	assign leaf[10949] = f[685] && f[239] && !f[322] && f[433];
	assign leaf[10950] = f[685] && f[239] && f[322] && !f[460];
	assign leaf[10951] = f[685] && f[239] && f[322] && f[460];
	
	// Tree 795, Classifier 5, Iteration: 79
	assign leaf[10952] = !f[411] && !f[468] && !f[354] && !f[301];
	assign leaf[10953] = !f[411] && !f[468] && !f[354] && f[301];
	assign leaf[10954] = !f[411] && !f[468] && f[354] && !f[324];
	assign leaf[10955] = !f[411] && !f[468] && f[354] && f[324];
	assign leaf[10956] = !f[411] && f[468] && !f[691] && !f[216];
	assign leaf[10957] = !f[411] && f[468] && !f[691] && f[216];
	assign leaf[10958] = !f[411] && f[468] && f[691];
	assign leaf[10959] = f[411] && !f[523] && !f[149] && !f[374];
	assign leaf[10960] = f[411] && !f[523] && !f[149] && f[374];
	assign leaf[10961] = f[411] && !f[523] && f[149] && !f[654];
	assign leaf[10962] = f[411] && !f[523] && f[149] && f[654];
	assign leaf[10963] = f[411] && f[523] && !f[187] && !f[157];
	assign leaf[10964] = f[411] && f[523] && !f[187] && f[157];
	assign leaf[10965] = f[411] && f[523] && f[187] && !f[237];
	assign leaf[10966] = f[411] && f[523] && f[187] && f[237];
	
	// Tree 796, Classifier 6, Iteration: 79
	assign leaf[10967] = !f[445] && !f[234] && !f[151] && !f[96];
	assign leaf[10968] = !f[445] && !f[234] && !f[151] && f[96];
	assign leaf[10969] = !f[445] && !f[234] && f[151] && !f[518];
	assign leaf[10970] = !f[445] && !f[234] && f[151] && f[518];
	assign leaf[10971] = !f[445] && f[234] && !f[373] && !f[426];
	assign leaf[10972] = !f[445] && f[234] && !f[373] && f[426];
	assign leaf[10973] = !f[445] && f[234] && f[373] && !f[152];
	assign leaf[10974] = !f[445] && f[234] && f[373] && f[152];
	assign leaf[10975] = f[445];
	
	// Tree 797, Classifier 7, Iteration: 79
	assign leaf[10976] = !f[437] && !f[273] && !f[176] && !f[517];
	assign leaf[10977] = !f[437] && !f[273] && !f[176] && f[517];
	assign leaf[10978] = !f[437] && !f[273] && f[176] && !f[494];
	assign leaf[10979] = !f[437] && !f[273] && f[176] && f[494];
	assign leaf[10980] = !f[437] && f[273] && !f[485] && !f[183];
	assign leaf[10981] = !f[437] && f[273] && !f[485] && f[183];
	assign leaf[10982] = !f[437] && f[273] && f[485];
	assign leaf[10983] = f[437] && !f[581] && !f[359] && !f[184];
	assign leaf[10984] = f[437] && !f[581] && !f[359] && f[184];
	assign leaf[10985] = f[437] && !f[581] && f[359] && !f[325];
	assign leaf[10986] = f[437] && !f[581] && f[359] && f[325];
	assign leaf[10987] = f[437] && f[581] && !f[204];
	assign leaf[10988] = f[437] && f[581] && f[204];
	
	// Tree 798, Classifier 8, Iteration: 79
	assign leaf[10989] = !f[317] && !f[518] && !f[295] && !f[321];
	assign leaf[10990] = !f[317] && !f[518] && !f[295] && f[321];
	assign leaf[10991] = !f[317] && !f[518] && f[295] && !f[236];
	assign leaf[10992] = !f[317] && !f[518] && f[295] && f[236];
	assign leaf[10993] = !f[317] && f[518] && !f[597] && !f[372];
	assign leaf[10994] = !f[317] && f[518] && !f[597] && f[372];
	assign leaf[10995] = !f[317] && f[518] && f[597] && !f[463];
	assign leaf[10996] = !f[317] && f[518] && f[597] && f[463];
	assign leaf[10997] = f[317] && !f[572] && !f[546] && !f[598];
	assign leaf[10998] = f[317] && !f[572] && !f[546] && f[598];
	assign leaf[10999] = f[317] && !f[572] && f[546] && !f[606];
	assign leaf[11000] = f[317] && !f[572] && f[546] && f[606];
	assign leaf[11001] = f[317] && f[572] && !f[685] && !f[431];
	assign leaf[11002] = f[317] && f[572] && !f[685] && f[431];
	assign leaf[11003] = f[317] && f[572] && f[685] && !f[580];
	assign leaf[11004] = f[317] && f[572] && f[685] && f[580];
	
	// Tree 799, Classifier 9, Iteration: 79
	assign leaf[11005] = !f[131] && !f[599] && !f[377] && !f[488];
	assign leaf[11006] = !f[131] && !f[599] && !f[377] && f[488];
	assign leaf[11007] = !f[131] && !f[599] && f[377] && !f[714];
	assign leaf[11008] = !f[131] && !f[599] && f[377] && f[714];
	assign leaf[11009] = !f[131] && f[599] && !f[487] && !f[378];
	assign leaf[11010] = !f[131] && f[599] && !f[487] && f[378];
	assign leaf[11011] = !f[131] && f[599] && f[487] && !f[434];
	assign leaf[11012] = !f[131] && f[599] && f[487] && f[434];
	assign leaf[11013] = f[131];
	
	// Tree 800, Classifier 0, Iteration: 80
	assign leaf[11014] = !f[526] && !f[635] && !f[688] && !f[378];
	assign leaf[11015] = !f[526] && !f[635] && !f[688] && f[378];
	assign leaf[11016] = !f[526] && !f[635] && f[688];
	assign leaf[11017] = !f[526] && f[635] && !f[578];
	assign leaf[11018] = !f[526] && f[635] && f[578] && !f[429];
	assign leaf[11019] = !f[526] && f[635] && f[578] && f[429];
	assign leaf[11020] = f[526] && !f[374] && !f[236] && !f[634];
	assign leaf[11021] = f[526] && !f[374] && !f[236] && f[634];
	assign leaf[11022] = f[526] && !f[374] && f[236] && !f[179];
	assign leaf[11023] = f[526] && !f[374] && f[236] && f[179];
	assign leaf[11024] = f[526] && f[374] && !f[544] && !f[233];
	assign leaf[11025] = f[526] && f[374] && !f[544] && f[233];
	assign leaf[11026] = f[526] && f[374] && f[544];
	
	// Tree 801, Classifier 1, Iteration: 80
	assign leaf[11027] = !f[440] && !f[204] && !f[658] && !f[517];
	assign leaf[11028] = !f[440] && !f[204] && !f[658] && f[517];
	assign leaf[11029] = !f[440] && !f[204] && f[658] && !f[436];
	assign leaf[11030] = !f[440] && !f[204] && f[658] && f[436];
	assign leaf[11031] = !f[440] && f[204] && !f[291] && !f[269];
	assign leaf[11032] = !f[440] && f[204] && !f[291] && f[269];
	assign leaf[11033] = !f[440] && f[204] && f[291];
	assign leaf[11034] = f[440];
	
	// Tree 802, Classifier 2, Iteration: 80
	assign leaf[11035] = !f[677] && !f[659] && !f[689] && !f[684];
	assign leaf[11036] = !f[677] && !f[659] && !f[689] && f[684];
	assign leaf[11037] = !f[677] && !f[659] && f[689] && !f[572];
	assign leaf[11038] = !f[677] && !f[659] && f[689] && f[572];
	assign leaf[11039] = !f[677] && f[659] && !f[465] && !f[269];
	assign leaf[11040] = !f[677] && f[659] && !f[465] && f[269];
	assign leaf[11041] = !f[677] && f[659] && f[465] && !f[229];
	assign leaf[11042] = !f[677] && f[659] && f[465] && f[229];
	assign leaf[11043] = f[677];
	
	// Tree 803, Classifier 3, Iteration: 80
	assign leaf[11044] = !f[209] && !f[265] && !f[261] && !f[235];
	assign leaf[11045] = !f[209] && !f[265] && !f[261] && f[235];
	assign leaf[11046] = !f[209] && !f[265] && f[261] && !f[470];
	assign leaf[11047] = !f[209] && !f[265] && f[261] && f[470];
	assign leaf[11048] = !f[209] && f[265] && !f[126] && !f[321];
	assign leaf[11049] = !f[209] && f[265] && !f[126] && f[321];
	assign leaf[11050] = !f[209] && f[265] && f[126] && !f[239];
	assign leaf[11051] = !f[209] && f[265] && f[126] && f[239];
	assign leaf[11052] = f[209] && !f[98] && !f[435] && !f[315];
	assign leaf[11053] = f[209] && !f[98] && !f[435] && f[315];
	assign leaf[11054] = f[209] && !f[98] && f[435] && !f[379];
	assign leaf[11055] = f[209] && !f[98] && f[435] && f[379];
	assign leaf[11056] = f[209] && f[98] && !f[123];
	assign leaf[11057] = f[209] && f[98] && f[123];
	
	// Tree 804, Classifier 4, Iteration: 80
	assign leaf[11058] = !f[385] && !f[320] && !f[237] && !f[181];
	assign leaf[11059] = !f[385] && !f[320] && !f[237] && f[181];
	assign leaf[11060] = !f[385] && !f[320] && f[237] && !f[154];
	assign leaf[11061] = !f[385] && !f[320] && f[237] && f[154];
	assign leaf[11062] = !f[385] && f[320] && !f[152] && !f[162];
	assign leaf[11063] = !f[385] && f[320] && !f[152] && f[162];
	assign leaf[11064] = !f[385] && f[320] && f[152] && !f[600];
	assign leaf[11065] = !f[385] && f[320] && f[152] && f[600];
	assign leaf[11066] = f[385] && !f[522] && !f[539] && !f[435];
	assign leaf[11067] = f[385] && !f[522] && !f[539] && f[435];
	assign leaf[11068] = f[385] && !f[522] && f[539] && !f[345];
	assign leaf[11069] = f[385] && !f[522] && f[539] && f[345];
	assign leaf[11070] = f[385] && f[522] && !f[353] && !f[464];
	assign leaf[11071] = f[385] && f[522] && !f[353] && f[464];
	assign leaf[11072] = f[385] && f[522] && f[353] && !f[518];
	assign leaf[11073] = f[385] && f[522] && f[353] && f[518];
	
	// Tree 805, Classifier 5, Iteration: 80
	assign leaf[11074] = !f[612] && !f[484] && !f[134] && !f[429];
	assign leaf[11075] = !f[612] && !f[484] && !f[134] && f[429];
	assign leaf[11076] = !f[612] && !f[484] && f[134] && !f[191];
	assign leaf[11077] = !f[612] && !f[484] && f[134] && f[191];
	assign leaf[11078] = !f[612] && f[484] && !f[429] && !f[459];
	assign leaf[11079] = !f[612] && f[484] && !f[429] && f[459];
	assign leaf[11080] = !f[612] && f[484] && f[429] && !f[540];
	assign leaf[11081] = !f[612] && f[484] && f[429] && f[540];
	assign leaf[11082] = f[612];
	
	// Tree 806, Classifier 6, Iteration: 80
	assign leaf[11083] = !f[517] && !f[234] && !f[151] && !f[242];
	assign leaf[11084] = !f[517] && !f[234] && !f[151] && f[242];
	assign leaf[11085] = !f[517] && !f[234] && f[151] && !f[347];
	assign leaf[11086] = !f[517] && !f[234] && f[151] && f[347];
	assign leaf[11087] = !f[517] && f[234] && !f[428] && !f[436];
	assign leaf[11088] = !f[517] && f[234] && !f[428] && f[436];
	assign leaf[11089] = !f[517] && f[234] && f[428] && !f[601];
	assign leaf[11090] = !f[517] && f[234] && f[428] && f[601];
	assign leaf[11091] = f[517] && !f[212] && !f[246] && !f[383];
	assign leaf[11092] = f[517] && !f[212] && !f[246] && f[383];
	assign leaf[11093] = f[517] && !f[212] && f[246] && !f[406];
	assign leaf[11094] = f[517] && !f[212] && f[246] && f[406];
	assign leaf[11095] = f[517] && f[212] && !f[599] && !f[551];
	assign leaf[11096] = f[517] && f[212] && !f[599] && f[551];
	assign leaf[11097] = f[517] && f[212] && f[599] && !f[521];
	assign leaf[11098] = f[517] && f[212] && f[599] && f[521];
	
	// Tree 807, Classifier 7, Iteration: 80
	assign leaf[11099] = !f[148] && !f[569] && !f[554] && !f[434];
	assign leaf[11100] = !f[148] && !f[569] && !f[554] && f[434];
	assign leaf[11101] = !f[148] && !f[569] && f[554] && !f[212];
	assign leaf[11102] = !f[148] && !f[569] && f[554] && f[212];
	assign leaf[11103] = !f[148] && f[569] && !f[651] && !f[260];
	assign leaf[11104] = !f[148] && f[569] && !f[651] && f[260];
	assign leaf[11105] = !f[148] && f[569] && f[651] && !f[547];
	assign leaf[11106] = !f[148] && f[569] && f[651] && f[547];
	assign leaf[11107] = f[148] && !f[324];
	assign leaf[11108] = f[148] && f[324] && !f[292] && !f[522];
	assign leaf[11109] = f[148] && f[324] && !f[292] && f[522];
	assign leaf[11110] = f[148] && f[324] && f[292];
	
	// Tree 808, Classifier 8, Iteration: 80
	assign leaf[11111] = !f[408] && !f[181] && !f[371] && !f[353];
	assign leaf[11112] = !f[408] && !f[181] && !f[371] && f[353];
	assign leaf[11113] = !f[408] && !f[181] && f[371] && !f[216];
	assign leaf[11114] = !f[408] && !f[181] && f[371] && f[216];
	assign leaf[11115] = !f[408] && f[181] && !f[268] && !f[158];
	assign leaf[11116] = !f[408] && f[181] && !f[268] && f[158];
	assign leaf[11117] = !f[408] && f[181] && f[268] && !f[602];
	assign leaf[11118] = !f[408] && f[181] && f[268] && f[602];
	assign leaf[11119] = f[408] && !f[577] && !f[324] && !f[465];
	assign leaf[11120] = f[408] && !f[577] && !f[324] && f[465];
	assign leaf[11121] = f[408] && !f[577] && f[324] && !f[435];
	assign leaf[11122] = f[408] && !f[577] && f[324] && f[435];
	assign leaf[11123] = f[408] && f[577] && !f[576] && !f[573];
	assign leaf[11124] = f[408] && f[577] && !f[576] && f[573];
	assign leaf[11125] = f[408] && f[577] && f[576] && !f[660];
	assign leaf[11126] = f[408] && f[577] && f[576] && f[660];
	
	// Tree 809, Classifier 9, Iteration: 80
	assign leaf[11127] = !f[244] && !f[275] && !f[327] && !f[213];
	assign leaf[11128] = !f[244] && !f[275] && !f[327] && f[213];
	assign leaf[11129] = !f[244] && !f[275] && f[327] && !f[211];
	assign leaf[11130] = !f[244] && !f[275] && f[327] && f[211];
	assign leaf[11131] = !f[244] && f[275] && !f[214];
	assign leaf[11132] = !f[244] && f[275] && f[214];
	assign leaf[11133] = f[244] && !f[385] && !f[209] && !f[299];
	assign leaf[11134] = f[244] && !f[385] && !f[209] && f[299];
	assign leaf[11135] = f[244] && !f[385] && f[209] && !f[185];
	assign leaf[11136] = f[244] && !f[385] && f[209] && f[185];
	assign leaf[11137] = f[244] && f[385] && !f[440] && !f[274];
	assign leaf[11138] = f[244] && f[385] && !f[440] && f[274];
	assign leaf[11139] = f[244] && f[385] && f[440] && !f[486];
	assign leaf[11140] = f[244] && f[385] && f[440] && f[486];
	
	// Tree 810, Classifier 0, Iteration: 81
	assign leaf[11141] = !f[386] && !f[497] && !f[354] && !f[511];
	assign leaf[11142] = !f[386] && !f[497] && !f[354] && f[511];
	assign leaf[11143] = !f[386] && !f[497] && f[354] && !f[509];
	assign leaf[11144] = !f[386] && !f[497] && f[354] && f[509];
	assign leaf[11145] = !f[386] && f[497] && !f[331] && !f[123];
	assign leaf[11146] = !f[386] && f[497] && !f[331] && f[123];
	assign leaf[11147] = !f[386] && f[497] && f[331];
	assign leaf[11148] = f[386] && !f[410] && !f[387] && !f[466];
	assign leaf[11149] = f[386] && !f[410] && !f[387] && f[466];
	assign leaf[11150] = f[386] && !f[410] && f[387] && !f[302];
	assign leaf[11151] = f[386] && !f[410] && f[387] && f[302];
	assign leaf[11152] = f[386] && f[410] && !f[513];
	assign leaf[11153] = f[386] && f[410] && f[513] && !f[297];
	assign leaf[11154] = f[386] && f[410] && f[513] && f[297];
	
	// Tree 811, Classifier 1, Iteration: 81
	assign leaf[11155] = !f[456] && !f[686] && !f[578] && !f[433];
	assign leaf[11156] = !f[456] && !f[686] && !f[578] && f[433];
	assign leaf[11157] = !f[456] && !f[686] && f[578] && !f[491];
	assign leaf[11158] = !f[456] && !f[686] && f[578] && f[491];
	assign leaf[11159] = !f[456] && f[686] && !f[180] && !f[263];
	assign leaf[11160] = !f[456] && f[686] && !f[180] && f[263];
	assign leaf[11161] = !f[456] && f[686] && f[180] && !f[347];
	assign leaf[11162] = !f[456] && f[686] && f[180] && f[347];
	assign leaf[11163] = f[456] && !f[630];
	assign leaf[11164] = f[456] && f[630];
	
	// Tree 812, Classifier 2, Iteration: 81
	assign leaf[11165] = !f[486] && !f[433] && !f[545] && !f[494];
	assign leaf[11166] = !f[486] && !f[433] && !f[545] && f[494];
	assign leaf[11167] = !f[486] && !f[433] && f[545] && !f[652];
	assign leaf[11168] = !f[486] && !f[433] && f[545] && f[652];
	assign leaf[11169] = !f[486] && f[433] && !f[456] && !f[491];
	assign leaf[11170] = !f[486] && f[433] && !f[456] && f[491];
	assign leaf[11171] = !f[486] && f[433] && f[456] && !f[325];
	assign leaf[11172] = !f[486] && f[433] && f[456] && f[325];
	assign leaf[11173] = f[486] && !f[432] && !f[324] && !f[568];
	assign leaf[11174] = f[486] && !f[432] && !f[324] && f[568];
	assign leaf[11175] = f[486] && !f[432] && f[324] && !f[601];
	assign leaf[11176] = f[486] && !f[432] && f[324] && f[601];
	assign leaf[11177] = f[486] && f[432] && !f[207] && !f[322];
	assign leaf[11178] = f[486] && f[432] && !f[207] && f[322];
	assign leaf[11179] = f[486] && f[432] && f[207] && !f[567];
	assign leaf[11180] = f[486] && f[432] && f[207] && f[567];
	
	// Tree 813, Classifier 3, Iteration: 81
	assign leaf[11181] = !f[429] && !f[96] && !f[178] && !f[241];
	assign leaf[11182] = !f[429] && !f[96] && !f[178] && f[241];
	assign leaf[11183] = !f[429] && !f[96] && f[178] && !f[261];
	assign leaf[11184] = !f[429] && !f[96] && f[178] && f[261];
	assign leaf[11185] = !f[429] && f[96] && !f[266] && !f[579];
	assign leaf[11186] = !f[429] && f[96] && !f[266] && f[579];
	assign leaf[11187] = !f[429] && f[96] && f[266] && !f[151];
	assign leaf[11188] = !f[429] && f[96] && f[266] && f[151];
	assign leaf[11189] = f[429] && !f[511] && !f[376] && !f[437];
	assign leaf[11190] = f[429] && !f[511] && !f[376] && f[437];
	assign leaf[11191] = f[429] && !f[511] && f[376] && !f[513];
	assign leaf[11192] = f[429] && !f[511] && f[376] && f[513];
	assign leaf[11193] = f[429] && f[511] && !f[542] && !f[434];
	assign leaf[11194] = f[429] && f[511] && !f[542] && f[434];
	assign leaf[11195] = f[429] && f[511] && f[542] && !f[181];
	assign leaf[11196] = f[429] && f[511] && f[542] && f[181];
	
	// Tree 814, Classifier 4, Iteration: 81
	assign leaf[11197] = !f[121] && !f[186] && !f[188] && !f[269];
	assign leaf[11198] = !f[121] && !f[186] && !f[188] && f[269];
	assign leaf[11199] = !f[121] && !f[186] && f[188] && !f[601];
	assign leaf[11200] = !f[121] && !f[186] && f[188] && f[601];
	assign leaf[11201] = !f[121] && f[186] && !f[269] && !f[295];
	assign leaf[11202] = !f[121] && f[186] && !f[269] && f[295];
	assign leaf[11203] = !f[121] && f[186] && f[269] && !f[469];
	assign leaf[11204] = !f[121] && f[186] && f[269] && f[469];
	assign leaf[11205] = f[121] && !f[574];
	assign leaf[11206] = f[121] && f[574];
	
	// Tree 815, Classifier 5, Iteration: 81
	assign leaf[11207] = !f[411] && !f[440] && !f[357] && !f[325];
	assign leaf[11208] = !f[411] && !f[440] && !f[357] && f[325];
	assign leaf[11209] = !f[411] && !f[440] && f[357] && !f[272];
	assign leaf[11210] = !f[411] && !f[440] && f[357] && f[272];
	assign leaf[11211] = !f[411] && f[440] && !f[635] && !f[319];
	assign leaf[11212] = !f[411] && f[440] && !f[635] && f[319];
	assign leaf[11213] = !f[411] && f[440] && f[635] && !f[210];
	assign leaf[11214] = !f[411] && f[440] && f[635] && f[210];
	assign leaf[11215] = f[411] && !f[329] && !f[185] && !f[127];
	assign leaf[11216] = f[411] && !f[329] && !f[185] && f[127];
	assign leaf[11217] = f[411] && !f[329] && f[185] && !f[271];
	assign leaf[11218] = f[411] && !f[329] && f[185] && f[271];
	assign leaf[11219] = f[411] && f[329] && !f[552];
	assign leaf[11220] = f[411] && f[329] && f[552];
	
	// Tree 816, Classifier 6, Iteration: 81
	assign leaf[11221] = !f[459] && !f[515] && !f[489] && !f[512];
	assign leaf[11222] = !f[459] && !f[515] && !f[489] && f[512];
	assign leaf[11223] = !f[459] && !f[515] && f[489] && !f[405];
	assign leaf[11224] = !f[459] && !f[515] && f[489] && f[405];
	assign leaf[11225] = !f[459] && f[515] && !f[359] && !f[457];
	assign leaf[11226] = !f[459] && f[515] && !f[359] && f[457];
	assign leaf[11227] = !f[459] && f[515] && f[359] && !f[407];
	assign leaf[11228] = !f[459] && f[515] && f[359] && f[407];
	assign leaf[11229] = f[459] && !f[610] && !f[316] && !f[687];
	assign leaf[11230] = f[459] && !f[610] && !f[316] && f[687];
	assign leaf[11231] = f[459] && !f[610] && f[316] && !f[384];
	assign leaf[11232] = f[459] && !f[610] && f[316] && f[384];
	assign leaf[11233] = f[459] && f[610];
	
	// Tree 817, Classifier 7, Iteration: 81
	assign leaf[11234] = !f[154] && !f[266] && !f[575] && !f[269];
	assign leaf[11235] = !f[154] && !f[266] && !f[575] && f[269];
	assign leaf[11236] = !f[154] && !f[266] && f[575] && !f[205];
	assign leaf[11237] = !f[154] && !f[266] && f[575] && f[205];
	assign leaf[11238] = !f[154] && f[266] && !f[263] && !f[294];
	assign leaf[11239] = !f[154] && f[266] && !f[263] && f[294];
	assign leaf[11240] = !f[154] && f[266] && f[263] && !f[368];
	assign leaf[11241] = !f[154] && f[266] && f[263] && f[368];
	assign leaf[11242] = f[154] && !f[463] && !f[571];
	assign leaf[11243] = f[154] && !f[463] && f[571];
	assign leaf[11244] = f[154] && f[463] && !f[403] && !f[236];
	assign leaf[11245] = f[154] && f[463] && !f[403] && f[236];
	assign leaf[11246] = f[154] && f[463] && f[403] && !f[152];
	assign leaf[11247] = f[154] && f[463] && f[403] && f[152];
	
	// Tree 818, Classifier 8, Iteration: 81
	assign leaf[11248] = !f[508] && !f[246] && !f[408] && !f[435];
	assign leaf[11249] = !f[508] && !f[246] && !f[408] && f[435];
	assign leaf[11250] = !f[508] && !f[246] && f[408] && !f[181];
	assign leaf[11251] = !f[508] && !f[246] && f[408] && f[181];
	assign leaf[11252] = !f[508] && f[246] && !f[329] && !f[215];
	assign leaf[11253] = !f[508] && f[246] && !f[329] && f[215];
	assign leaf[11254] = !f[508] && f[246] && f[329] && !f[374];
	assign leaf[11255] = !f[508] && f[246] && f[329] && f[374];
	assign leaf[11256] = f[508] && !f[153];
	assign leaf[11257] = f[508] && f[153];
	
	// Tree 819, Classifier 9, Iteration: 81
	assign leaf[11258] = !f[201] && !f[632] && !f[128] && !f[292];
	assign leaf[11259] = !f[201] && !f[632] && !f[128] && f[292];
	assign leaf[11260] = !f[201] && !f[632] && f[128];
	assign leaf[11261] = !f[201] && f[632] && !f[546] && !f[155];
	assign leaf[11262] = !f[201] && f[632] && !f[546] && f[155];
	assign leaf[11263] = !f[201] && f[632] && f[546] && !f[513];
	assign leaf[11264] = !f[201] && f[632] && f[546] && f[513];
	assign leaf[11265] = f[201] && !f[428];
	assign leaf[11266] = f[201] && f[428];
	
	// Tree 820, Classifier 0, Iteration: 82
	assign leaf[11267] = !f[434] && !f[459] && !f[349] && !f[547];
	assign leaf[11268] = !f[434] && !f[459] && !f[349] && f[547];
	assign leaf[11269] = !f[434] && !f[459] && f[349] && !f[426];
	assign leaf[11270] = !f[434] && !f[459] && f[349] && f[426];
	assign leaf[11271] = !f[434] && f[459] && !f[601] && !f[484];
	assign leaf[11272] = !f[434] && f[459] && !f[601] && f[484];
	assign leaf[11273] = !f[434] && f[459] && f[601] && !f[656];
	assign leaf[11274] = !f[434] && f[459] && f[601] && f[656];
	assign leaf[11275] = f[434] && !f[433];
	assign leaf[11276] = f[434] && f[433] && !f[431];
	assign leaf[11277] = f[434] && f[433] && f[431] && !f[521];
	assign leaf[11278] = f[434] && f[433] && f[431] && f[521];
	
	// Tree 821, Classifier 1, Iteration: 82
	assign leaf[11279] = !f[329] && !f[375] && !f[321] && !f[181];
	assign leaf[11280] = !f[329] && !f[375] && !f[321] && f[181];
	assign leaf[11281] = !f[329] && !f[375] && f[321] && !f[622];
	assign leaf[11282] = !f[329] && !f[375] && f[321] && f[622];
	assign leaf[11283] = !f[329] && f[375] && !f[321] && !f[548];
	assign leaf[11284] = !f[329] && f[375] && !f[321] && f[548];
	assign leaf[11285] = !f[329] && f[375] && f[321] && !f[658];
	assign leaf[11286] = !f[329] && f[375] && f[321] && f[658];
	assign leaf[11287] = f[329];
	
	// Tree 822, Classifier 2, Iteration: 82
	assign leaf[11288] = !f[121] && !f[528] && !f[500] && !f[388];
	assign leaf[11289] = !f[121] && !f[528] && !f[500] && f[388];
	assign leaf[11290] = !f[121] && !f[528] && f[500] && !f[241];
	assign leaf[11291] = !f[121] && !f[528] && f[500] && f[241];
	assign leaf[11292] = !f[121] && f[528] && !f[500] && !f[512];
	assign leaf[11293] = !f[121] && f[528] && !f[500] && f[512];
	assign leaf[11294] = !f[121] && f[528] && f[500] && !f[319];
	assign leaf[11295] = !f[121] && f[528] && f[500] && f[319];
	assign leaf[11296] = f[121] && !f[289] && !f[633] && !f[605];
	assign leaf[11297] = f[121] && !f[289] && !f[633] && f[605];
	assign leaf[11298] = f[121] && !f[289] && f[633] && !f[498];
	assign leaf[11299] = f[121] && !f[289] && f[633] && f[498];
	assign leaf[11300] = f[121] && f[289];
	
	// Tree 823, Classifier 3, Iteration: 82
	assign leaf[11301] = !f[705] && !f[358] && !f[330] && !f[357];
	assign leaf[11302] = !f[705] && !f[358] && !f[330] && f[357];
	assign leaf[11303] = !f[705] && !f[358] && f[330] && !f[321];
	assign leaf[11304] = !f[705] && !f[358] && f[330] && f[321];
	assign leaf[11305] = !f[705] && f[358] && !f[595];
	assign leaf[11306] = !f[705] && f[358] && f[595] && !f[576];
	assign leaf[11307] = !f[705] && f[358] && f[595] && f[576];
	assign leaf[11308] = f[705];
	
	// Tree 824, Classifier 4, Iteration: 82
	assign leaf[11309] = !f[738] && !f[72] && !f[94] && !f[383];
	assign leaf[11310] = !f[738] && !f[72] && !f[94] && f[383];
	assign leaf[11311] = !f[738] && !f[72] && f[94];
	assign leaf[11312] = !f[738] && f[72];
	assign leaf[11313] = f[738];
	
	// Tree 825, Classifier 5, Iteration: 82
	assign leaf[11314] = !f[402] && !f[187] && !f[239] && !f[128];
	assign leaf[11315] = !f[402] && !f[187] && !f[239] && f[128];
	assign leaf[11316] = !f[402] && !f[187] && f[239] && !f[244];
	assign leaf[11317] = !f[402] && !f[187] && f[239] && f[244];
	assign leaf[11318] = !f[402] && f[187] && !f[211] && !f[215];
	assign leaf[11319] = !f[402] && f[187] && !f[211] && f[215];
	assign leaf[11320] = !f[402] && f[187] && f[211] && !f[299];
	assign leaf[11321] = !f[402] && f[187] && f[211] && f[299];
	assign leaf[11322] = f[402] && !f[484] && !f[568] && !f[491];
	assign leaf[11323] = f[402] && !f[484] && !f[568] && f[491];
	assign leaf[11324] = f[402] && !f[484] && f[568] && !f[319];
	assign leaf[11325] = f[402] && !f[484] && f[568] && f[319];
	assign leaf[11326] = f[402] && f[484] && !f[625] && !f[638];
	assign leaf[11327] = f[402] && f[484] && !f[625] && f[638];
	assign leaf[11328] = f[402] && f[484] && f[625] && !f[467];
	assign leaf[11329] = f[402] && f[484] && f[625] && f[467];
	
	// Tree 826, Classifier 6, Iteration: 82
	assign leaf[11330] = !f[652] && !f[267] && !f[237] && !f[183];
	assign leaf[11331] = !f[652] && !f[267] && !f[237] && f[183];
	assign leaf[11332] = !f[652] && !f[267] && f[237] && !f[328];
	assign leaf[11333] = !f[652] && !f[267] && f[237] && f[328];
	assign leaf[11334] = !f[652] && f[267] && !f[321] && !f[545];
	assign leaf[11335] = !f[652] && f[267] && !f[321] && f[545];
	assign leaf[11336] = !f[652] && f[267] && f[321] && !f[580];
	assign leaf[11337] = !f[652] && f[267] && f[321] && f[580];
	assign leaf[11338] = f[652] && !f[512];
	assign leaf[11339] = f[652] && f[512];
	
	// Tree 827, Classifier 7, Iteration: 82
	assign leaf[11340] = !f[686] && !f[575] && !f[683] && !f[518];
	assign leaf[11341] = !f[686] && !f[575] && !f[683] && f[518];
	assign leaf[11342] = !f[686] && !f[575] && f[683] && !f[624];
	assign leaf[11343] = !f[686] && !f[575] && f[683] && f[624];
	assign leaf[11344] = !f[686] && f[575] && !f[492] && !f[203];
	assign leaf[11345] = !f[686] && f[575] && !f[492] && f[203];
	assign leaf[11346] = !f[686] && f[575] && f[492] && !f[259];
	assign leaf[11347] = !f[686] && f[575] && f[492] && f[259];
	assign leaf[11348] = f[686] && !f[682] && !f[661] && !f[323];
	assign leaf[11349] = f[686] && !f[682] && !f[661] && f[323];
	assign leaf[11350] = f[686] && !f[682] && f[661] && !f[716];
	assign leaf[11351] = f[686] && !f[682] && f[661] && f[716];
	assign leaf[11352] = f[686] && f[682] && !f[301] && !f[573];
	assign leaf[11353] = f[686] && f[682] && !f[301] && f[573];
	assign leaf[11354] = f[686] && f[682] && f[301];
	
	// Tree 828, Classifier 8, Iteration: 82
	assign leaf[11355] = !f[302] && !f[235] && !f[234] && !f[348];
	assign leaf[11356] = !f[302] && !f[235] && !f[234] && f[348];
	assign leaf[11357] = !f[302] && !f[235] && f[234] && !f[291];
	assign leaf[11358] = !f[302] && !f[235] && f[234] && f[291];
	assign leaf[11359] = !f[302] && f[235] && !f[320] && !f[375];
	assign leaf[11360] = !f[302] && f[235] && !f[320] && f[375];
	assign leaf[11361] = !f[302] && f[235] && f[320] && !f[349];
	assign leaf[11362] = !f[302] && f[235] && f[320] && f[349];
	assign leaf[11363] = f[302] && !f[457] && !f[402] && !f[377];
	assign leaf[11364] = f[302] && !f[457] && !f[402] && f[377];
	assign leaf[11365] = f[302] && !f[457] && f[402] && !f[404];
	assign leaf[11366] = f[302] && !f[457] && f[402] && f[404];
	assign leaf[11367] = f[302] && f[457] && !f[443] && !f[329];
	assign leaf[11368] = f[302] && f[457] && !f[443] && f[329];
	assign leaf[11369] = f[302] && f[457] && f[443];
	
	// Tree 829, Classifier 9, Iteration: 82
	assign leaf[11370] = !f[599] && !f[543] && !f[540] && !f[740];
	assign leaf[11371] = !f[599] && !f[543] && !f[540] && f[740];
	assign leaf[11372] = !f[599] && !f[543] && f[540] && !f[482];
	assign leaf[11373] = !f[599] && !f[543] && f[540] && f[482];
	assign leaf[11374] = !f[599] && f[543] && !f[432] && !f[459];
	assign leaf[11375] = !f[599] && f[543] && !f[432] && f[459];
	assign leaf[11376] = !f[599] && f[543] && f[432] && !f[428];
	assign leaf[11377] = !f[599] && f[543] && f[432] && f[428];
	assign leaf[11378] = f[599] && !f[488] && !f[272] && !f[511];
	assign leaf[11379] = f[599] && !f[488] && !f[272] && f[511];
	assign leaf[11380] = f[599] && !f[488] && f[272] && !f[238];
	assign leaf[11381] = f[599] && !f[488] && f[272] && f[238];
	assign leaf[11382] = f[599] && f[488] && !f[186] && !f[516];
	assign leaf[11383] = f[599] && f[488] && !f[186] && f[516];
	assign leaf[11384] = f[599] && f[488] && f[186] && !f[680];
	assign leaf[11385] = f[599] && f[488] && f[186] && f[680];
	
	// Tree 830, Classifier 0, Iteration: 83
	assign leaf[11386] = !f[380] && !f[512] && !f[629] && !f[290];
	assign leaf[11387] = !f[380] && !f[512] && !f[629] && f[290];
	assign leaf[11388] = !f[380] && !f[512] && f[629] && !f[209];
	assign leaf[11389] = !f[380] && !f[512] && f[629] && f[209];
	assign leaf[11390] = !f[380] && f[512] && !f[302] && !f[517];
	assign leaf[11391] = !f[380] && f[512] && !f[302] && f[517];
	assign leaf[11392] = !f[380] && f[512] && f[302] && !f[271];
	assign leaf[11393] = !f[380] && f[512] && f[302] && f[271];
	assign leaf[11394] = f[380] && !f[297] && !f[184];
	assign leaf[11395] = f[380] && !f[297] && f[184];
	assign leaf[11396] = f[380] && f[297] && !f[435] && !f[262];
	assign leaf[11397] = f[380] && f[297] && !f[435] && f[262];
	assign leaf[11398] = f[380] && f[297] && f[435] && !f[406];
	assign leaf[11399] = f[380] && f[297] && f[435] && f[406];
	
	// Tree 831, Classifier 1, Iteration: 83
	assign leaf[11400] = !f[709] && !f[204] && !f[245] && !f[538];
	assign leaf[11401] = !f[709] && !f[204] && !f[245] && f[538];
	assign leaf[11402] = !f[709] && !f[204] && f[245] && !f[162];
	assign leaf[11403] = !f[709] && !f[204] && f[245] && f[162];
	assign leaf[11404] = !f[709] && f[204] && !f[569] && !f[636];
	assign leaf[11405] = !f[709] && f[204] && !f[569] && f[636];
	assign leaf[11406] = !f[709] && f[204] && f[569];
	assign leaf[11407] = f[709];
	
	// Tree 832, Classifier 2, Iteration: 83
	assign leaf[11408] = !f[154] && !f[99] && !f[377] && !f[372];
	assign leaf[11409] = !f[154] && !f[99] && !f[377] && f[372];
	assign leaf[11410] = !f[154] && !f[99] && f[377] && !f[484];
	assign leaf[11411] = !f[154] && !f[99] && f[377] && f[484];
	assign leaf[11412] = !f[154] && f[99] && !f[566] && !f[487];
	assign leaf[11413] = !f[154] && f[99] && !f[566] && f[487];
	assign leaf[11414] = !f[154] && f[99] && f[566];
	assign leaf[11415] = f[154] && !f[636] && !f[294] && !f[625];
	assign leaf[11416] = f[154] && !f[636] && !f[294] && f[625];
	assign leaf[11417] = f[154] && !f[636] && f[294] && !f[553];
	assign leaf[11418] = f[154] && !f[636] && f[294] && f[553];
	assign leaf[11419] = f[154] && f[636] && !f[524] && !f[526];
	assign leaf[11420] = f[154] && f[636] && !f[524] && f[526];
	assign leaf[11421] = f[154] && f[636] && f[524] && !f[662];
	assign leaf[11422] = f[154] && f[636] && f[524] && f[662];
	
	// Tree 833, Classifier 3, Iteration: 83
	assign leaf[11423] = !f[377] && !f[324] && !f[436] && !f[321];
	assign leaf[11424] = !f[377] && !f[324] && !f[436] && f[321];
	assign leaf[11425] = !f[377] && !f[324] && f[436] && !f[539];
	assign leaf[11426] = !f[377] && !f[324] && f[436] && f[539];
	assign leaf[11427] = !f[377] && f[324] && !f[436] && !f[547];
	assign leaf[11428] = !f[377] && f[324] && !f[436] && f[547];
	assign leaf[11429] = !f[377] && f[324] && f[436] && !f[604];
	assign leaf[11430] = !f[377] && f[324] && f[436] && f[604];
	assign leaf[11431] = f[377] && !f[181] && !f[126] && !f[263];
	assign leaf[11432] = f[377] && !f[181] && !f[126] && f[263];
	assign leaf[11433] = f[377] && !f[181] && f[126] && !f[436];
	assign leaf[11434] = f[377] && !f[181] && f[126] && f[436];
	assign leaf[11435] = f[377] && f[181] && !f[264] && !f[290];
	assign leaf[11436] = f[377] && f[181] && !f[264] && f[290];
	assign leaf[11437] = f[377] && f[181] && f[264] && !f[316];
	assign leaf[11438] = f[377] && f[181] && f[264] && f[316];
	
	// Tree 834, Classifier 4, Iteration: 83
	assign leaf[11439] = !f[384] && !f[494] && !f[435] && !f[294];
	assign leaf[11440] = !f[384] && !f[494] && !f[435] && f[294];
	assign leaf[11441] = !f[384] && !f[494] && f[435] && !f[326];
	assign leaf[11442] = !f[384] && !f[494] && f[435] && f[326];
	assign leaf[11443] = !f[384] && f[494] && !f[206] && !f[518];
	assign leaf[11444] = !f[384] && f[494] && !f[206] && f[518];
	assign leaf[11445] = !f[384] && f[494] && f[206] && !f[210];
	assign leaf[11446] = !f[384] && f[494] && f[206] && f[210];
	assign leaf[11447] = f[384] && !f[439] && !f[486] && !f[351];
	assign leaf[11448] = f[384] && !f[439] && !f[486] && f[351];
	assign leaf[11449] = f[384] && !f[439] && f[486] && !f[210];
	assign leaf[11450] = f[384] && !f[439] && f[486] && f[210];
	assign leaf[11451] = f[384] && f[439] && !f[353] && !f[214];
	assign leaf[11452] = f[384] && f[439] && !f[353] && f[214];
	assign leaf[11453] = f[384] && f[439] && f[353] && !f[271];
	assign leaf[11454] = f[384] && f[439] && f[353] && f[271];
	
	// Tree 835, Classifier 5, Iteration: 83
	assign leaf[11455] = !f[276] && !f[380] && !f[681] && !f[521];
	assign leaf[11456] = !f[276] && !f[380] && !f[681] && f[521];
	assign leaf[11457] = !f[276] && !f[380] && f[681] && !f[548];
	assign leaf[11458] = !f[276] && !f[380] && f[681] && f[548];
	assign leaf[11459] = !f[276] && f[380] && !f[328] && !f[131];
	assign leaf[11460] = !f[276] && f[380] && !f[328] && f[131];
	assign leaf[11461] = !f[276] && f[380] && f[328] && !f[407];
	assign leaf[11462] = !f[276] && f[380] && f[328] && f[407];
	assign leaf[11463] = f[276] && !f[273];
	assign leaf[11464] = f[276] && f[273] && !f[234] && !f[351];
	assign leaf[11465] = f[276] && f[273] && !f[234] && f[351];
	assign leaf[11466] = f[276] && f[273] && f[234];
	
	// Tree 836, Classifier 6, Iteration: 83
	assign leaf[11467] = !f[299] && !f[301] && !f[272] && !f[383];
	assign leaf[11468] = !f[299] && !f[301] && !f[272] && f[383];
	assign leaf[11469] = !f[299] && !f[301] && f[272];
	assign leaf[11470] = !f[299] && f[301] && !f[403] && !f[434];
	assign leaf[11471] = !f[299] && f[301] && !f[403] && f[434];
	assign leaf[11472] = !f[299] && f[301] && f[403];
	assign leaf[11473] = f[299] && !f[382] && !f[658] && !f[388];
	assign leaf[11474] = f[299] && !f[382] && !f[658] && f[388];
	assign leaf[11475] = f[299] && !f[382] && f[658] && !f[293];
	assign leaf[11476] = f[299] && !f[382] && f[658] && f[293];
	assign leaf[11477] = f[299] && f[382] && !f[352] && !f[301];
	assign leaf[11478] = f[299] && f[382] && !f[352] && f[301];
	assign leaf[11479] = f[299] && f[382] && f[352] && !f[494];
	assign leaf[11480] = f[299] && f[382] && f[352] && f[494];
	
	// Tree 837, Classifier 7, Iteration: 83
	assign leaf[11481] = !f[238] && !f[235] && !f[322] && !f[208];
	assign leaf[11482] = !f[238] && !f[235] && !f[322] && f[208];
	assign leaf[11483] = !f[238] && !f[235] && f[322] && !f[318];
	assign leaf[11484] = !f[238] && !f[235] && f[322] && f[318];
	assign leaf[11485] = !f[238] && f[235] && !f[208] && !f[436];
	assign leaf[11486] = !f[238] && f[235] && !f[208] && f[436];
	assign leaf[11487] = !f[238] && f[235] && f[208] && !f[546];
	assign leaf[11488] = !f[238] && f[235] && f[208] && f[546];
	assign leaf[11489] = f[238] && !f[236] && !f[718] && !f[401];
	assign leaf[11490] = f[238] && !f[236] && !f[718] && f[401];
	assign leaf[11491] = f[238] && !f[236] && f[718];
	assign leaf[11492] = f[238] && f[236] && !f[329] && !f[214];
	assign leaf[11493] = f[238] && f[236] && !f[329] && f[214];
	assign leaf[11494] = f[238] && f[236] && f[329] && !f[274];
	assign leaf[11495] = f[238] && f[236] && f[329] && f[274];
	
	// Tree 838, Classifier 8, Iteration: 83
	assign leaf[11496] = !f[469] && !f[386] && !f[453] && !f[133];
	assign leaf[11497] = !f[469] && !f[386] && !f[453] && f[133];
	assign leaf[11498] = !f[469] && !f[386] && f[453];
	assign leaf[11499] = !f[469] && f[386] && !f[375] && !f[577];
	assign leaf[11500] = !f[469] && f[386] && !f[375] && f[577];
	assign leaf[11501] = !f[469] && f[386] && f[375] && !f[300];
	assign leaf[11502] = !f[469] && f[386] && f[375] && f[300];
	assign leaf[11503] = f[469] && !f[523] && !f[299] && !f[459];
	assign leaf[11504] = f[469] && !f[523] && !f[299] && f[459];
	assign leaf[11505] = f[469] && !f[523] && f[299] && !f[411];
	assign leaf[11506] = f[469] && !f[523] && f[299] && f[411];
	assign leaf[11507] = f[469] && f[523] && !f[183] && !f[151];
	assign leaf[11508] = f[469] && f[523] && !f[183] && f[151];
	assign leaf[11509] = f[469] && f[523] && f[183] && !f[593];
	assign leaf[11510] = f[469] && f[523] && f[183] && f[593];
	
	// Tree 839, Classifier 9, Iteration: 83
	assign leaf[11511] = !f[744] && !f[524] && !f[469] && !f[379];
	assign leaf[11512] = !f[744] && !f[524] && !f[469] && f[379];
	assign leaf[11513] = !f[744] && !f[524] && f[469] && !f[413];
	assign leaf[11514] = !f[744] && !f[524] && f[469] && f[413];
	assign leaf[11515] = !f[744] && f[524] && !f[259] && !f[565];
	assign leaf[11516] = !f[744] && f[524] && !f[259] && f[565];
	assign leaf[11517] = !f[744] && f[524] && f[259] && !f[290];
	assign leaf[11518] = !f[744] && f[524] && f[259] && f[290];
	assign leaf[11519] = f[744] && !f[434] && !f[322] && !f[351];
	assign leaf[11520] = f[744] && !f[434] && !f[322] && f[351];
	assign leaf[11521] = f[744] && !f[434] && f[322];
	assign leaf[11522] = f[744] && f[434] && !f[690] && !f[287];
	assign leaf[11523] = f[744] && f[434] && !f[690] && f[287];
	assign leaf[11524] = f[744] && f[434] && f[690];
	
	// Tree 840, Classifier 0, Iteration: 84
	assign leaf[11525] = !f[152] && !f[294] && !f[155] && !f[488];
	assign leaf[11526] = !f[152] && !f[294] && !f[155] && f[488];
	assign leaf[11527] = !f[152] && !f[294] && f[155] && !f[463];
	assign leaf[11528] = !f[152] && !f[294] && f[155] && f[463];
	assign leaf[11529] = !f[152] && f[294] && !f[100] && !f[351];
	assign leaf[11530] = !f[152] && f[294] && !f[100] && f[351];
	assign leaf[11531] = !f[152] && f[294] && f[100];
	assign leaf[11532] = f[152] && !f[371] && !f[539] && !f[156];
	assign leaf[11533] = f[152] && !f[371] && !f[539] && f[156];
	assign leaf[11534] = f[152] && !f[371] && f[539] && !f[465];
	assign leaf[11535] = f[152] && !f[371] && f[539] && f[465];
	assign leaf[11536] = f[152] && f[371] && !f[455];
	assign leaf[11537] = f[152] && f[371] && f[455] && !f[214];
	assign leaf[11538] = f[152] && f[371] && f[455] && f[214];
	
	// Tree 841, Classifier 1, Iteration: 84
	assign leaf[11539] = !f[708] && !f[244] && !f[204] && !f[266];
	assign leaf[11540] = !f[708] && !f[244] && !f[204] && f[266];
	assign leaf[11541] = !f[708] && !f[244] && f[204] && !f[156];
	assign leaf[11542] = !f[708] && !f[244] && f[204] && f[156];
	assign leaf[11543] = !f[708] && f[244] && !f[293] && !f[129];
	assign leaf[11544] = !f[708] && f[244] && !f[293] && f[129];
	assign leaf[11545] = !f[708] && f[244] && f[293] && !f[595];
	assign leaf[11546] = !f[708] && f[244] && f[293] && f[595];
	assign leaf[11547] = f[708];
	
	// Tree 842, Classifier 2, Iteration: 84
	assign leaf[11548] = !f[417] && !f[351] && !f[355] && !f[228];
	assign leaf[11549] = !f[417] && !f[351] && !f[355] && f[228];
	assign leaf[11550] = !f[417] && !f[351] && f[355] && !f[384];
	assign leaf[11551] = !f[417] && !f[351] && f[355] && f[384];
	assign leaf[11552] = !f[417] && f[351] && !f[606] && !f[216];
	assign leaf[11553] = !f[417] && f[351] && !f[606] && f[216];
	assign leaf[11554] = !f[417] && f[351] && f[606] && !f[205];
	assign leaf[11555] = !f[417] && f[351] && f[606] && f[205];
	assign leaf[11556] = f[417] && !f[240];
	assign leaf[11557] = f[417] && f[240];
	
	// Tree 843, Classifier 3, Iteration: 84
	assign leaf[11558] = !f[315] && !f[259] && !f[150] && !f[325];
	assign leaf[11559] = !f[315] && !f[259] && !f[150] && f[325];
	assign leaf[11560] = !f[315] && !f[259] && f[150] && !f[233];
	assign leaf[11561] = !f[315] && !f[259] && f[150] && f[233];
	assign leaf[11562] = !f[315] && f[259] && !f[375] && !f[572];
	assign leaf[11563] = !f[315] && f[259] && !f[375] && f[572];
	assign leaf[11564] = !f[315] && f[259] && f[375] && !f[149];
	assign leaf[11565] = !f[315] && f[259] && f[375] && f[149];
	assign leaf[11566] = f[315] && !f[345] && !f[399] && !f[433];
	assign leaf[11567] = f[315] && !f[345] && !f[399] && f[433];
	assign leaf[11568] = f[315] && !f[345] && f[399];
	assign leaf[11569] = f[315] && f[345] && !f[291] && !f[625];
	assign leaf[11570] = f[315] && f[345] && !f[291] && f[625];
	assign leaf[11571] = f[315] && f[345] && f[291] && !f[238];
	assign leaf[11572] = f[315] && f[345] && f[291] && f[238];
	
	// Tree 844, Classifier 4, Iteration: 84
	assign leaf[11573] = !f[275] && !f[123] && !f[238] && !f[240];
	assign leaf[11574] = !f[275] && !f[123] && !f[238] && f[240];
	assign leaf[11575] = !f[275] && !f[123] && f[238] && !f[154];
	assign leaf[11576] = !f[275] && !f[123] && f[238] && f[154];
	assign leaf[11577] = !f[275] && f[123] && !f[484];
	assign leaf[11578] = !f[275] && f[123] && f[484];
	assign leaf[11579] = f[275] && !f[453] && !f[385] && !f[237];
	assign leaf[11580] = f[275] && !f[453] && !f[385] && f[237];
	assign leaf[11581] = f[275] && !f[453] && f[385] && !f[245];
	assign leaf[11582] = f[275] && !f[453] && f[385] && f[245];
	assign leaf[11583] = f[275] && f[453];
	
	// Tree 845, Classifier 5, Iteration: 84
	assign leaf[11584] = !f[216] && !f[322] && !f[599] && !f[524];
	assign leaf[11585] = !f[216] && !f[322] && !f[599] && f[524];
	assign leaf[11586] = !f[216] && !f[322] && f[599] && !f[242];
	assign leaf[11587] = !f[216] && !f[322] && f[599] && f[242];
	assign leaf[11588] = !f[216] && f[322] && !f[267] && !f[242];
	assign leaf[11589] = !f[216] && f[322] && !f[267] && f[242];
	assign leaf[11590] = !f[216] && f[322] && f[267] && !f[299];
	assign leaf[11591] = !f[216] && f[322] && f[267] && f[299];
	assign leaf[11592] = f[216] && !f[299] && !f[370] && !f[213];
	assign leaf[11593] = f[216] && !f[299] && !f[370] && f[213];
	assign leaf[11594] = f[216] && !f[299] && f[370] && !f[662];
	assign leaf[11595] = f[216] && !f[299] && f[370] && f[662];
	assign leaf[11596] = f[216] && f[299] && !f[268];
	assign leaf[11597] = f[216] && f[299] && f[268] && !f[272];
	assign leaf[11598] = f[216] && f[299] && f[268] && f[272];
	
	// Tree 846, Classifier 6, Iteration: 84
	assign leaf[11599] = !f[571] && !f[575] && !f[399] && !f[187];
	assign leaf[11600] = !f[571] && !f[575] && !f[399] && f[187];
	assign leaf[11601] = !f[571] && !f[575] && f[399] && !f[401];
	assign leaf[11602] = !f[571] && !f[575] && f[399] && f[401];
	assign leaf[11603] = !f[571] && f[575] && !f[659] && !f[242];
	assign leaf[11604] = !f[571] && f[575] && !f[659] && f[242];
	assign leaf[11605] = !f[571] && f[575] && f[659] && !f[545];
	assign leaf[11606] = !f[571] && f[575] && f[659] && f[545];
	assign leaf[11607] = f[571] && !f[486] && !f[181] && !f[98];
	assign leaf[11608] = f[571] && !f[486] && !f[181] && f[98];
	assign leaf[11609] = f[571] && !f[486] && f[181] && !f[315];
	assign leaf[11610] = f[571] && !f[486] && f[181] && f[315];
	assign leaf[11611] = f[571] && f[486] && !f[687] && !f[568];
	assign leaf[11612] = f[571] && f[486] && !f[687] && f[568];
	assign leaf[11613] = f[571] && f[486] && f[687];
	
	// Tree 847, Classifier 7, Iteration: 84
	assign leaf[11614] = !f[464] && !f[574] && !f[300] && !f[236];
	assign leaf[11615] = !f[464] && !f[574] && !f[300] && f[236];
	assign leaf[11616] = !f[464] && !f[574] && f[300] && !f[683];
	assign leaf[11617] = !f[464] && !f[574] && f[300] && f[683];
	assign leaf[11618] = !f[464] && f[574] && !f[377] && !f[492];
	assign leaf[11619] = !f[464] && f[574] && !f[377] && f[492];
	assign leaf[11620] = !f[464] && f[574] && f[377] && !f[659];
	assign leaf[11621] = !f[464] && f[574] && f[377] && f[659];
	assign leaf[11622] = f[464] && !f[595] && !f[518] && !f[682];
	assign leaf[11623] = f[464] && !f[595] && !f[518] && f[682];
	assign leaf[11624] = f[464] && !f[595] && f[518] && !f[269];
	assign leaf[11625] = f[464] && !f[595] && f[518] && f[269];
	assign leaf[11626] = f[464] && f[595] && !f[677] && !f[440];
	assign leaf[11627] = f[464] && f[595] && !f[677] && f[440];
	assign leaf[11628] = f[464] && f[595] && f[677];
	
	// Tree 848, Classifier 8, Iteration: 84
	assign leaf[11629] = !f[525] && !f[629] && !f[684] && !f[608];
	assign leaf[11630] = !f[525] && !f[629] && !f[684] && f[608];
	assign leaf[11631] = !f[525] && !f[629] && f[684] && !f[464];
	assign leaf[11632] = !f[525] && !f[629] && f[684] && f[464];
	assign leaf[11633] = !f[525] && f[629] && !f[657] && !f[572];
	assign leaf[11634] = !f[525] && f[629] && !f[657] && f[572];
	assign leaf[11635] = !f[525] && f[629] && f[657] && !f[543];
	assign leaf[11636] = !f[525] && f[629] && f[657] && f[543];
	assign leaf[11637] = f[525] && !f[458] && !f[571] && !f[522];
	assign leaf[11638] = f[525] && !f[458] && !f[571] && f[522];
	assign leaf[11639] = f[525] && !f[458] && f[571] && !f[689];
	assign leaf[11640] = f[525] && !f[458] && f[571] && f[689];
	assign leaf[11641] = f[525] && f[458] && !f[322] && !f[624];
	assign leaf[11642] = f[525] && f[458] && !f[322] && f[624];
	assign leaf[11643] = f[525] && f[458] && f[322] && !f[385];
	assign leaf[11644] = f[525] && f[458] && f[322] && f[385];
	
	// Tree 849, Classifier 9, Iteration: 84
	assign leaf[11645] = !f[508] && !f[350] && !f[340] && !f[401];
	assign leaf[11646] = !f[508] && !f[350] && !f[340] && f[401];
	assign leaf[11647] = !f[508] && !f[350] && f[340] && !f[212];
	assign leaf[11648] = !f[508] && !f[350] && f[340] && f[212];
	assign leaf[11649] = !f[508] && f[350] && !f[352] && !f[267];
	assign leaf[11650] = !f[508] && f[350] && !f[352] && f[267];
	assign leaf[11651] = !f[508] && f[350] && f[352] && !f[402];
	assign leaf[11652] = !f[508] && f[350] && f[352] && f[402];
	assign leaf[11653] = f[508];
	
	// Tree 850, Classifier 0, Iteration: 85
	assign leaf[11654] = !f[681] && !f[345] && !f[375] && !f[498];
	assign leaf[11655] = !f[681] && !f[345] && !f[375] && f[498];
	assign leaf[11656] = !f[681] && !f[345] && f[375] && !f[429];
	assign leaf[11657] = !f[681] && !f[345] && f[375] && f[429];
	assign leaf[11658] = !f[681] && f[345] && !f[376] && !f[570];
	assign leaf[11659] = !f[681] && f[345] && !f[376] && f[570];
	assign leaf[11660] = !f[681] && f[345] && f[376] && !f[264];
	assign leaf[11661] = !f[681] && f[345] && f[376] && f[264];
	assign leaf[11662] = f[681] && !f[599] && !f[354] && !f[523];
	assign leaf[11663] = f[681] && !f[599] && !f[354] && f[523];
	assign leaf[11664] = f[681] && !f[599] && f[354];
	assign leaf[11665] = f[681] && f[599] && !f[575];
	assign leaf[11666] = f[681] && f[599] && f[575];
	
	// Tree 851, Classifier 1, Iteration: 85
	assign leaf[11667] = !f[493] && !f[519] && !f[464] && !f[353];
	assign leaf[11668] = !f[493] && !f[519] && !f[464] && f[353];
	assign leaf[11669] = !f[493] && !f[519] && f[464] && !f[487];
	assign leaf[11670] = !f[493] && !f[519] && f[464] && f[487];
	assign leaf[11671] = !f[493] && f[519] && !f[546] && !f[180];
	assign leaf[11672] = !f[493] && f[519] && !f[546] && f[180];
	assign leaf[11673] = !f[493] && f[519] && f[546] && !f[462];
	assign leaf[11674] = !f[493] && f[519] && f[546] && f[462];
	assign leaf[11675] = f[493] && !f[636] && !f[547];
	assign leaf[11676] = f[493] && !f[636] && f[547] && !f[265];
	assign leaf[11677] = f[493] && !f[636] && f[547] && f[265];
	assign leaf[11678] = f[493] && f[636];
	
	// Tree 852, Classifier 2, Iteration: 85
	assign leaf[11679] = !f[709] && !f[712] && !f[134] && !f[104];
	assign leaf[11680] = !f[709] && !f[712] && !f[134] && f[104];
	assign leaf[11681] = !f[709] && !f[712] && f[134] && !f[273];
	assign leaf[11682] = !f[709] && !f[712] && f[134] && f[273];
	assign leaf[11683] = !f[709] && f[712];
	assign leaf[11684] = f[709];
	
	// Tree 853, Classifier 3, Iteration: 85
	assign leaf[11685] = !f[406] && !f[315] && !f[517] && !f[348];
	assign leaf[11686] = !f[406] && !f[315] && !f[517] && f[348];
	assign leaf[11687] = !f[406] && !f[315] && f[517] && !f[296];
	assign leaf[11688] = !f[406] && !f[315] && f[517] && f[296];
	assign leaf[11689] = !f[406] && f[315] && !f[438] && !f[327];
	assign leaf[11690] = !f[406] && f[315] && !f[438] && f[327];
	assign leaf[11691] = !f[406] && f[315] && f[438] && !f[489];
	assign leaf[11692] = !f[406] && f[315] && f[438] && f[489];
	assign leaf[11693] = f[406] && !f[604] && !f[608] && !f[547];
	assign leaf[11694] = f[406] && !f[604] && !f[608] && f[547];
	assign leaf[11695] = f[406] && !f[604] && f[608] && !f[235];
	assign leaf[11696] = f[406] && !f[604] && f[608] && f[235];
	assign leaf[11697] = f[406] && f[604] && !f[346] && !f[380];
	assign leaf[11698] = f[406] && f[604] && !f[346] && f[380];
	assign leaf[11699] = f[406] && f[604] && f[346] && !f[403];
	assign leaf[11700] = f[406] && f[604] && f[346] && f[403];
	
	// Tree 854, Classifier 4, Iteration: 85
	assign leaf[11701] = !f[663] && !f[606] && !f[579] && !f[513];
	assign leaf[11702] = !f[663] && !f[606] && !f[579] && f[513];
	assign leaf[11703] = !f[663] && !f[606] && f[579] && !f[213];
	assign leaf[11704] = !f[663] && !f[606] && f[579] && f[213];
	assign leaf[11705] = !f[663] && f[606] && !f[549];
	assign leaf[11706] = !f[663] && f[606] && f[549] && !f[349];
	assign leaf[11707] = !f[663] && f[606] && f[549] && f[349];
	assign leaf[11708] = f[663] && !f[462] && !f[267] && !f[578];
	assign leaf[11709] = f[663] && !f[462] && !f[267] && f[578];
	assign leaf[11710] = f[663] && !f[462] && f[267] && !f[464];
	assign leaf[11711] = f[663] && !f[462] && f[267] && f[464];
	assign leaf[11712] = f[663] && f[462] && !f[206] && !f[290];
	assign leaf[11713] = f[663] && f[462] && !f[206] && f[290];
	assign leaf[11714] = f[663] && f[462] && f[206] && !f[232];
	assign leaf[11715] = f[663] && f[462] && f[206] && f[232];
	
	// Tree 855, Classifier 5, Iteration: 85
	assign leaf[11716] = !f[717] && !f[577] && !f[432] && !f[411];
	assign leaf[11717] = !f[717] && !f[577] && !f[432] && f[411];
	assign leaf[11718] = !f[717] && !f[577] && f[432] && !f[330];
	assign leaf[11719] = !f[717] && !f[577] && f[432] && f[330];
	assign leaf[11720] = !f[717] && f[577] && !f[397] && !f[216];
	assign leaf[11721] = !f[717] && f[577] && !f[397] && f[216];
	assign leaf[11722] = !f[717] && f[577] && f[397] && !f[353];
	assign leaf[11723] = !f[717] && f[577] && f[397] && f[353];
	assign leaf[11724] = f[717] && !f[351] && !f[577];
	assign leaf[11725] = f[717] && !f[351] && f[577];
	assign leaf[11726] = f[717] && f[351];
	
	// Tree 856, Classifier 6, Iteration: 85
	assign leaf[11727] = !f[247] && !f[574] && !f[570] && !f[571];
	assign leaf[11728] = !f[247] && !f[574] && !f[570] && f[571];
	assign leaf[11729] = !f[247] && !f[574] && f[570] && !f[152];
	assign leaf[11730] = !f[247] && !f[574] && f[570] && f[152];
	assign leaf[11731] = !f[247] && f[574] && !f[209] && !f[320];
	assign leaf[11732] = !f[247] && f[574] && !f[209] && f[320];
	assign leaf[11733] = !f[247] && f[574] && f[209] && !f[126];
	assign leaf[11734] = !f[247] && f[574] && f[209] && f[126];
	assign leaf[11735] = f[247] && !f[630];
	assign leaf[11736] = f[247] && f[630];
	
	// Tree 857, Classifier 7, Iteration: 85
	assign leaf[11737] = !f[510] && !f[609] && !f[291] && !f[288];
	assign leaf[11738] = !f[510] && !f[609] && !f[291] && f[288];
	assign leaf[11739] = !f[510] && !f[609] && f[291] && !f[287];
	assign leaf[11740] = !f[510] && !f[609] && f[291] && f[287];
	assign leaf[11741] = !f[510] && f[609] && !f[349];
	assign leaf[11742] = !f[510] && f[609] && f[349];
	assign leaf[11743] = f[510] && !f[685] && !f[342] && !f[267];
	assign leaf[11744] = f[510] && !f[685] && !f[342] && f[267];
	assign leaf[11745] = f[510] && !f[685] && f[342];
	assign leaf[11746] = f[510] && f[685];
	
	// Tree 858, Classifier 8, Iteration: 85
	assign leaf[11747] = !f[214] && !f[434] && !f[379] && !f[435];
	assign leaf[11748] = !f[214] && !f[434] && !f[379] && f[435];
	assign leaf[11749] = !f[214] && !f[434] && f[379] && !f[271];
	assign leaf[11750] = !f[214] && !f[434] && f[379] && f[271];
	assign leaf[11751] = !f[214] && f[434] && !f[293] && !f[348];
	assign leaf[11752] = !f[214] && f[434] && !f[293] && f[348];
	assign leaf[11753] = !f[214] && f[434] && f[293] && !f[187];
	assign leaf[11754] = !f[214] && f[434] && f[293] && f[187];
	assign leaf[11755] = f[214] && !f[212] && !f[211] && !f[188];
	assign leaf[11756] = f[214] && !f[212] && !f[211] && f[188];
	assign leaf[11757] = f[214] && !f[212] && f[211] && !f[239];
	assign leaf[11758] = f[214] && !f[212] && f[211] && f[239];
	assign leaf[11759] = f[214] && f[212] && !f[329] && !f[482];
	assign leaf[11760] = f[214] && f[212] && !f[329] && f[482];
	assign leaf[11761] = f[214] && f[212] && f[329] && !f[273];
	assign leaf[11762] = f[214] && f[212] && f[329] && f[273];
	
	// Tree 859, Classifier 9, Iteration: 85
	assign leaf[11763] = !f[742] && !f[407] && !f[346] && !f[574];
	assign leaf[11764] = !f[742] && !f[407] && !f[346] && f[574];
	assign leaf[11765] = !f[742] && !f[407] && f[346] && !f[432];
	assign leaf[11766] = !f[742] && !f[407] && f[346] && f[432];
	assign leaf[11767] = !f[742] && f[407] && !f[291] && !f[211];
	assign leaf[11768] = !f[742] && f[407] && !f[291] && f[211];
	assign leaf[11769] = !f[742] && f[407] && f[291] && !f[206];
	assign leaf[11770] = !f[742] && f[407] && f[291] && f[206];
	assign leaf[11771] = f[742] && !f[573] && !f[315] && !f[379];
	assign leaf[11772] = f[742] && !f[573] && !f[315] && f[379];
	assign leaf[11773] = f[742] && !f[573] && f[315] && !f[209];
	assign leaf[11774] = f[742] && !f[573] && f[315] && f[209];
	assign leaf[11775] = f[742] && f[573] && !f[458];
	assign leaf[11776] = f[742] && f[573] && f[458];
	
	// Tree 860, Classifier 0, Iteration: 86
	assign leaf[11777] = !f[633] && !f[683] && !f[608] && !f[378];
	assign leaf[11778] = !f[633] && !f[683] && !f[608] && f[378];
	assign leaf[11779] = !f[633] && !f[683] && f[608];
	assign leaf[11780] = !f[633] && f[683] && !f[156];
	assign leaf[11781] = !f[633] && f[683] && f[156] && !f[235];
	assign leaf[11782] = !f[633] && f[683] && f[156] && f[235];
	assign leaf[11783] = f[633] && !f[579] && !f[576];
	assign leaf[11784] = f[633] && !f[579] && f[576] && !f[542];
	assign leaf[11785] = f[633] && !f[579] && f[576] && f[542];
	assign leaf[11786] = f[633] && f[579] && !f[234] && !f[266];
	assign leaf[11787] = f[633] && f[579] && !f[234] && f[266];
	assign leaf[11788] = f[633] && f[579] && f[234] && !f[157];
	assign leaf[11789] = f[633] && f[579] && f[234] && f[157];
	
	// Tree 861, Classifier 1, Iteration: 86
	assign leaf[11790] = !f[356] && !f[215] && !f[353] && !f[566];
	assign leaf[11791] = !f[356] && !f[215] && !f[353] && f[566];
	assign leaf[11792] = !f[356] && !f[215] && f[353] && !f[659];
	assign leaf[11793] = !f[356] && !f[215] && f[353] && f[659];
	assign leaf[11794] = !f[356] && f[215] && !f[381] && !f[519];
	assign leaf[11795] = !f[356] && f[215] && !f[381] && f[519];
	assign leaf[11796] = !f[356] && f[215] && f[381] && !f[436];
	assign leaf[11797] = !f[356] && f[215] && f[381] && f[436];
	assign leaf[11798] = f[356];
	
	// Tree 862, Classifier 2, Iteration: 86
	assign leaf[11799] = !f[374] && !f[125] && !f[209] && !f[326];
	assign leaf[11800] = !f[374] && !f[125] && !f[209] && f[326];
	assign leaf[11801] = !f[374] && !f[125] && f[209] && !f[599];
	assign leaf[11802] = !f[374] && !f[125] && f[209] && f[599];
	assign leaf[11803] = !f[374] && f[125] && !f[594] && !f[213];
	assign leaf[11804] = !f[374] && f[125] && !f[594] && f[213];
	assign leaf[11805] = !f[374] && f[125] && f[594] && !f[578];
	assign leaf[11806] = !f[374] && f[125] && f[594] && f[578];
	assign leaf[11807] = f[374] && !f[398] && !f[127] && !f[470];
	assign leaf[11808] = f[374] && !f[398] && !f[127] && f[470];
	assign leaf[11809] = f[374] && !f[398] && f[127] && !f[129];
	assign leaf[11810] = f[374] && !f[398] && f[127] && f[129];
	assign leaf[11811] = f[374] && f[398] && !f[323] && !f[573];
	assign leaf[11812] = f[374] && f[398] && !f[323] && f[573];
	assign leaf[11813] = f[374] && f[398] && f[323];
	
	// Tree 863, Classifier 3, Iteration: 86
	assign leaf[11814] = !f[386] && !f[401] && !f[347] && !f[290];
	assign leaf[11815] = !f[386] && !f[401] && !f[347] && f[290];
	assign leaf[11816] = !f[386] && !f[401] && f[347] && !f[459];
	assign leaf[11817] = !f[386] && !f[401] && f[347] && f[459];
	assign leaf[11818] = !f[386] && f[401] && !f[509] && !f[442];
	assign leaf[11819] = !f[386] && f[401] && !f[509] && f[442];
	assign leaf[11820] = !f[386] && f[401] && f[509] && !f[454];
	assign leaf[11821] = !f[386] && f[401] && f[509] && f[454];
	assign leaf[11822] = f[386] && !f[499];
	assign leaf[11823] = f[386] && f[499] && !f[287];
	assign leaf[11824] = f[386] && f[499] && f[287];
	
	// Tree 864, Classifier 4, Iteration: 86
	assign leaf[11825] = !f[184] && !f[182] && !f[294] && !f[239];
	assign leaf[11826] = !f[184] && !f[182] && !f[294] && f[239];
	assign leaf[11827] = !f[184] && !f[182] && f[294] && !f[291];
	assign leaf[11828] = !f[184] && !f[182] && f[294] && f[291];
	assign leaf[11829] = !f[184] && f[182] && !f[206] && !f[294];
	assign leaf[11830] = !f[184] && f[182] && !f[206] && f[294];
	assign leaf[11831] = !f[184] && f[182] && f[206] && !f[291];
	assign leaf[11832] = !f[184] && f[182] && f[206] && f[291];
	assign leaf[11833] = f[184] && !f[215] && !f[239] && !f[268];
	assign leaf[11834] = f[184] && !f[215] && !f[239] && f[268];
	assign leaf[11835] = f[184] && !f[215] && f[239] && !f[159];
	assign leaf[11836] = f[184] && !f[215] && f[239] && f[159];
	assign leaf[11837] = f[184] && f[215] && !f[581] && !f[441];
	assign leaf[11838] = f[184] && f[215] && !f[581] && f[441];
	assign leaf[11839] = f[184] && f[215] && f[581];
	
	// Tree 865, Classifier 5, Iteration: 86
	assign leaf[11840] = !f[685] && !f[521] && !f[205] && !f[318];
	assign leaf[11841] = !f[685] && !f[521] && !f[205] && f[318];
	assign leaf[11842] = !f[685] && !f[521] && f[205] && !f[375];
	assign leaf[11843] = !f[685] && !f[521] && f[205] && f[375];
	assign leaf[11844] = !f[685] && f[521] && !f[234] && !f[548];
	assign leaf[11845] = !f[685] && f[521] && !f[234] && f[548];
	assign leaf[11846] = !f[685] && f[521] && f[234] && !f[127];
	assign leaf[11847] = !f[685] && f[521] && f[234] && f[127];
	assign leaf[11848] = f[685] && !f[546] && !f[290] && !f[294];
	assign leaf[11849] = f[685] && !f[546] && !f[290] && f[294];
	assign leaf[11850] = f[685] && !f[546] && f[290] && !f[174];
	assign leaf[11851] = f[685] && !f[546] && f[290] && f[174];
	assign leaf[11852] = f[685] && f[546] && !f[210];
	assign leaf[11853] = f[685] && f[546] && f[210] && !f[274];
	assign leaf[11854] = f[685] && f[546] && f[210] && f[274];
	
	// Tree 866, Classifier 6, Iteration: 86
	assign leaf[11855] = !f[107] && !f[214] && !f[293] && !f[155];
	assign leaf[11856] = !f[107] && !f[214] && !f[293] && f[155];
	assign leaf[11857] = !f[107] && !f[214] && f[293] && !f[156];
	assign leaf[11858] = !f[107] && !f[214] && f[293] && f[156];
	assign leaf[11859] = !f[107] && f[214] && !f[433] && !f[509];
	assign leaf[11860] = !f[107] && f[214] && !f[433] && f[509];
	assign leaf[11861] = !f[107] && f[214] && f[433] && !f[352];
	assign leaf[11862] = !f[107] && f[214] && f[433] && f[352];
	assign leaf[11863] = f[107];
	
	// Tree 867, Classifier 7, Iteration: 86
	assign leaf[11864] = !f[707] && !f[625] && !f[600] && !f[682];
	assign leaf[11865] = !f[707] && !f[625] && !f[600] && f[682];
	assign leaf[11866] = !f[707] && !f[625] && f[600] && !f[318];
	assign leaf[11867] = !f[707] && !f[625] && f[600] && f[318];
	assign leaf[11868] = !f[707] && f[625] && !f[602] && !f[685];
	assign leaf[11869] = !f[707] && f[625] && !f[602] && f[685];
	assign leaf[11870] = !f[707] && f[625] && f[602] && !f[685];
	assign leaf[11871] = !f[707] && f[625] && f[602] && f[685];
	assign leaf[11872] = f[707] && !f[597] && !f[706] && !f[185];
	assign leaf[11873] = f[707] && !f[597] && !f[706] && f[185];
	assign leaf[11874] = f[707] && !f[597] && f[706];
	assign leaf[11875] = f[707] && f[597] && !f[348] && !f[318];
	assign leaf[11876] = f[707] && f[597] && !f[348] && f[318];
	assign leaf[11877] = f[707] && f[597] && f[348];
	
	// Tree 868, Classifier 8, Iteration: 86
	assign leaf[11878] = !f[125] && !f[439] && !f[525] && !f[592];
	assign leaf[11879] = !f[125] && !f[439] && !f[525] && f[592];
	assign leaf[11880] = !f[125] && !f[439] && f[525] && !f[187];
	assign leaf[11881] = !f[125] && !f[439] && f[525] && f[187];
	assign leaf[11882] = !f[125] && f[439] && !f[521] && !f[324];
	assign leaf[11883] = !f[125] && f[439] && !f[521] && f[324];
	assign leaf[11884] = !f[125] && f[439] && f[521] && !f[303];
	assign leaf[11885] = !f[125] && f[439] && f[521] && f[303];
	assign leaf[11886] = f[125] && !f[128] && !f[273] && !f[378];
	assign leaf[11887] = f[125] && !f[128] && !f[273] && f[378];
	assign leaf[11888] = f[125] && !f[128] && f[273];
	assign leaf[11889] = f[125] && f[128] && !f[431] && !f[605];
	assign leaf[11890] = f[125] && f[128] && !f[431] && f[605];
	assign leaf[11891] = f[125] && f[128] && f[431] && !f[296];
	assign leaf[11892] = f[125] && f[128] && f[431] && f[296];
	
	// Tree 869, Classifier 9, Iteration: 86
	assign leaf[11893] = !f[500] && !f[162] && !f[122] && !f[686];
	assign leaf[11894] = !f[500] && !f[162] && !f[122] && f[686];
	assign leaf[11895] = !f[500] && !f[162] && f[122];
	assign leaf[11896] = !f[500] && f[162];
	assign leaf[11897] = f[500];
	
	// Tree 870, Classifier 0, Iteration: 87
	assign leaf[11898] = !f[380] && !f[456] && !f[516] && !f[212];
	assign leaf[11899] = !f[380] && !f[456] && !f[516] && f[212];
	assign leaf[11900] = !f[380] && !f[456] && f[516] && !f[266];
	assign leaf[11901] = !f[380] && !f[456] && f[516] && f[266];
	assign leaf[11902] = !f[380] && f[456] && !f[654] && !f[520];
	assign leaf[11903] = !f[380] && f[456] && !f[654] && f[520];
	assign leaf[11904] = !f[380] && f[456] && f[654] && !f[681];
	assign leaf[11905] = !f[380] && f[456] && f[654] && f[681];
	assign leaf[11906] = f[380] && !f[378] && !f[377] && !f[412];
	assign leaf[11907] = f[380] && !f[378] && !f[377] && f[412];
	assign leaf[11908] = f[380] && !f[378] && f[377];
	assign leaf[11909] = f[380] && f[378] && !f[427] && !f[410];
	assign leaf[11910] = f[380] && f[378] && !f[427] && f[410];
	assign leaf[11911] = f[380] && f[378] && f[427] && !f[273];
	assign leaf[11912] = f[380] && f[378] && f[427] && f[273];
	
	// Tree 871, Classifier 1, Iteration: 87
	assign leaf[11913] = !f[152] && !f[656] && !f[573] && !f[714];
	assign leaf[11914] = !f[152] && !f[656] && !f[573] && f[714];
	assign leaf[11915] = !f[152] && !f[656] && f[573] && !f[486];
	assign leaf[11916] = !f[152] && !f[656] && f[573] && f[486];
	assign leaf[11917] = !f[152] && f[656] && !f[380] && !f[270];
	assign leaf[11918] = !f[152] && f[656] && !f[380] && f[270];
	assign leaf[11919] = !f[152] && f[656] && f[380] && !f[463];
	assign leaf[11920] = !f[152] && f[656] && f[380] && f[463];
	assign leaf[11921] = f[152] && !f[269] && !f[236] && !f[206];
	assign leaf[11922] = f[152] && !f[269] && !f[236] && f[206];
	assign leaf[11923] = f[152] && !f[269] && f[236] && !f[547];
	assign leaf[11924] = f[152] && !f[269] && f[236] && f[547];
	assign leaf[11925] = f[152] && f[269] && !f[462];
	assign leaf[11926] = f[152] && f[269] && f[462] && !f[375];
	assign leaf[11927] = f[152] && f[269] && f[462] && f[375];
	
	// Tree 872, Classifier 2, Iteration: 87
	assign leaf[11928] = !f[413] && !f[572] && !f[322] && !f[233];
	assign leaf[11929] = !f[413] && !f[572] && !f[322] && f[233];
	assign leaf[11930] = !f[413] && !f[572] && f[322] && !f[525];
	assign leaf[11931] = !f[413] && !f[572] && f[322] && f[525];
	assign leaf[11932] = !f[413] && f[572] && !f[406] && !f[540];
	assign leaf[11933] = !f[413] && f[572] && !f[406] && f[540];
	assign leaf[11934] = !f[413] && f[572] && f[406] && !f[681];
	assign leaf[11935] = !f[413] && f[572] && f[406] && f[681];
	assign leaf[11936] = f[413] && !f[464] && !f[174] && !f[624];
	assign leaf[11937] = f[413] && !f[464] && !f[174] && f[624];
	assign leaf[11938] = f[413] && !f[464] && f[174];
	assign leaf[11939] = f[413] && f[464] && !f[490] && !f[212];
	assign leaf[11940] = f[413] && f[464] && !f[490] && f[212];
	assign leaf[11941] = f[413] && f[464] && f[490] && !f[242];
	assign leaf[11942] = f[413] && f[464] && f[490] && f[242];
	
	// Tree 873, Classifier 3, Iteration: 87
	assign leaf[11943] = !f[707] && !f[344] && !f[270] && !f[187];
	assign leaf[11944] = !f[707] && !f[344] && !f[270] && f[187];
	assign leaf[11945] = !f[707] && !f[344] && f[270] && !f[293];
	assign leaf[11946] = !f[707] && !f[344] && f[270] && f[293];
	assign leaf[11947] = !f[707] && f[344] && !f[402] && !f[636];
	assign leaf[11948] = !f[707] && f[344] && !f[402] && f[636];
	assign leaf[11949] = !f[707] && f[344] && f[402] && !f[347];
	assign leaf[11950] = !f[707] && f[344] && f[402] && f[347];
	assign leaf[11951] = f[707] && !f[267];
	assign leaf[11952] = f[707] && f[267] && !f[493];
	assign leaf[11953] = f[707] && f[267] && f[493];
	
	// Tree 874, Classifier 4, Iteration: 87
	assign leaf[11954] = !f[746] && !f[429] && !f[349] && !f[188];
	assign leaf[11955] = !f[746] && !f[429] && !f[349] && f[188];
	assign leaf[11956] = !f[746] && !f[429] && f[349] && !f[466];
	assign leaf[11957] = !f[746] && !f[429] && f[349] && f[466];
	assign leaf[11958] = !f[746] && f[429] && !f[397] && !f[374];
	assign leaf[11959] = !f[746] && f[429] && !f[397] && f[374];
	assign leaf[11960] = !f[746] && f[429] && f[397] && !f[382];
	assign leaf[11961] = !f[746] && f[429] && f[397] && f[382];
	assign leaf[11962] = f[746];
	
	// Tree 875, Classifier 5, Iteration: 87
	assign leaf[11963] = !f[333] && !f[622] && !f[598] && !f[654];
	assign leaf[11964] = !f[333] && !f[622] && !f[598] && f[654];
	assign leaf[11965] = !f[333] && !f[622] && f[598] && !f[397];
	assign leaf[11966] = !f[333] && !f[622] && f[598] && f[397];
	assign leaf[11967] = !f[333] && f[622] && !f[540] && !f[179];
	assign leaf[11968] = !f[333] && f[622] && !f[540] && f[179];
	assign leaf[11969] = !f[333] && f[622] && f[540] && !f[537];
	assign leaf[11970] = !f[333] && f[622] && f[540] && f[537];
	assign leaf[11971] = f[333];
	
	// Tree 876, Classifier 6, Iteration: 87
	assign leaf[11972] = !f[299] && !f[301] && !f[383] && !f[123];
	assign leaf[11973] = !f[299] && !f[301] && !f[383] && f[123];
	assign leaf[11974] = !f[299] && !f[301] && f[383] && !f[405];
	assign leaf[11975] = !f[299] && !f[301] && f[383] && f[405];
	assign leaf[11976] = !f[299] && f[301] && !f[489];
	assign leaf[11977] = !f[299] && f[301] && f[489] && !f[289];
	assign leaf[11978] = !f[299] && f[301] && f[489] && f[289];
	assign leaf[11979] = f[299] && !f[358] && !f[348] && !f[233];
	assign leaf[11980] = f[299] && !f[358] && !f[348] && f[233];
	assign leaf[11981] = f[299] && !f[358] && f[348] && !f[542];
	assign leaf[11982] = f[299] && !f[358] && f[348] && f[542];
	assign leaf[11983] = f[299] && f[358] && !f[600];
	assign leaf[11984] = f[299] && f[358] && f[600] && !f[486];
	assign leaf[11985] = f[299] && f[358] && f[600] && f[486];
	
	// Tree 877, Classifier 7, Iteration: 87
	assign leaf[11986] = !f[434] && !f[488] && !f[458] && !f[432];
	assign leaf[11987] = !f[434] && !f[488] && !f[458] && f[432];
	assign leaf[11988] = !f[434] && !f[488] && f[458] && !f[374];
	assign leaf[11989] = !f[434] && !f[488] && f[458] && f[374];
	assign leaf[11990] = !f[434] && f[488] && !f[430] && !f[412];
	assign leaf[11991] = !f[434] && f[488] && !f[430] && f[412];
	assign leaf[11992] = !f[434] && f[488] && f[430] && !f[494];
	assign leaf[11993] = !f[434] && f[488] && f[430] && f[494];
	assign leaf[11994] = f[434] && !f[606] && !f[320] && !f[346];
	assign leaf[11995] = f[434] && !f[606] && !f[320] && f[346];
	assign leaf[11996] = f[434] && !f[606] && f[320] && !f[210];
	assign leaf[11997] = f[434] && !f[606] && f[320] && f[210];
	assign leaf[11998] = f[434] && f[606] && !f[202];
	assign leaf[11999] = f[434] && f[606] && f[202] && !f[327];
	assign leaf[12000] = f[434] && f[606] && f[202] && f[327];
	
	// Tree 878, Classifier 8, Iteration: 87
	assign leaf[12001] = !f[692] && !f[689] && !f[688] && !f[715];
	assign leaf[12002] = !f[692] && !f[689] && !f[688] && f[715];
	assign leaf[12003] = !f[692] && !f[689] && f[688] && !f[631];
	assign leaf[12004] = !f[692] && !f[689] && f[688] && f[631];
	assign leaf[12005] = !f[692] && f[689] && !f[493] && !f[631];
	assign leaf[12006] = !f[692] && f[689] && !f[493] && f[631];
	assign leaf[12007] = !f[692] && f[689] && f[493] && !f[272];
	assign leaf[12008] = !f[692] && f[689] && f[493] && f[272];
	assign leaf[12009] = f[692] && !f[268] && !f[238];
	assign leaf[12010] = f[692] && !f[268] && f[238];
	assign leaf[12011] = f[692] && f[268] && !f[575] && !f[460];
	assign leaf[12012] = f[692] && f[268] && !f[575] && f[460];
	assign leaf[12013] = f[692] && f[268] && f[575];
	
	// Tree 879, Classifier 9, Iteration: 87
	assign leaf[12014] = !f[742] && !f[351] && !f[433] && !f[489];
	assign leaf[12015] = !f[742] && !f[351] && !f[433] && f[489];
	assign leaf[12016] = !f[742] && !f[351] && f[433] && !f[516];
	assign leaf[12017] = !f[742] && !f[351] && f[433] && f[516];
	assign leaf[12018] = !f[742] && f[351] && !f[353] && !f[409];
	assign leaf[12019] = !f[742] && f[351] && !f[353] && f[409];
	assign leaf[12020] = !f[742] && f[351] && f[353] && !f[385];
	assign leaf[12021] = !f[742] && f[351] && f[353] && f[385];
	assign leaf[12022] = f[742] && !f[290] && !f[407];
	assign leaf[12023] = f[742] && !f[290] && f[407] && !f[294];
	assign leaf[12024] = f[742] && !f[290] && f[407] && f[294];
	assign leaf[12025] = f[742] && f[290] && !f[234] && !f[399];
	assign leaf[12026] = f[742] && f[290] && !f[234] && f[399];
	assign leaf[12027] = f[742] && f[290] && f[234] && !f[461];
	assign leaf[12028] = f[742] && f[290] && f[234] && f[461];
	
	// Tree 880, Classifier 0, Iteration: 88
	assign leaf[12029] = !f[514] && !f[539] && !f[513] && !f[508];
	assign leaf[12030] = !f[514] && !f[539] && !f[513] && f[508];
	assign leaf[12031] = !f[514] && !f[539] && f[513] && !f[185];
	assign leaf[12032] = !f[514] && !f[539] && f[513] && f[185];
	assign leaf[12033] = !f[514] && f[539] && !f[624] && !f[183];
	assign leaf[12034] = !f[514] && f[539] && !f[624] && f[183];
	assign leaf[12035] = !f[514] && f[539] && f[624] && !f[483];
	assign leaf[12036] = !f[514] && f[539] && f[624] && f[483];
	assign leaf[12037] = f[514] && !f[567] && !f[465] && !f[349];
	assign leaf[12038] = f[514] && !f[567] && !f[465] && f[349];
	assign leaf[12039] = f[514] && !f[567] && f[465] && !f[268];
	assign leaf[12040] = f[514] && !f[567] && f[465] && f[268];
	assign leaf[12041] = f[514] && f[567] && !f[371] && !f[651];
	assign leaf[12042] = f[514] && f[567] && !f[371] && f[651];
	assign leaf[12043] = f[514] && f[567] && f[371];
	
	// Tree 881, Classifier 1, Iteration: 88
	assign leaf[12044] = !f[244] && !f[566] && !f[493] && !f[178];
	assign leaf[12045] = !f[244] && !f[566] && !f[493] && f[178];
	assign leaf[12046] = !f[244] && !f[566] && f[493] && !f[519];
	assign leaf[12047] = !f[244] && !f[566] && f[493] && f[519];
	assign leaf[12048] = !f[244] && f[566] && !f[349];
	assign leaf[12049] = !f[244] && f[566] && f[349];
	assign leaf[12050] = f[244] && !f[321] && !f[381];
	assign leaf[12051] = f[244] && !f[321] && f[381] && !f[296];
	assign leaf[12052] = f[244] && !f[321] && f[381] && f[296];
	assign leaf[12053] = f[244] && f[321] && !f[320] && !f[430];
	assign leaf[12054] = f[244] && f[321] && !f[320] && f[430];
	assign leaf[12055] = f[244] && f[321] && f[320];
	
	// Tree 882, Classifier 2, Iteration: 88
	assign leaf[12056] = !f[486] && !f[432] && !f[209] && !f[492];
	assign leaf[12057] = !f[486] && !f[432] && !f[209] && f[492];
	assign leaf[12058] = !f[486] && !f[432] && f[209] && !f[568];
	assign leaf[12059] = !f[486] && !f[432] && f[209] && f[568];
	assign leaf[12060] = !f[486] && f[432] && !f[456] && !f[436];
	assign leaf[12061] = !f[486] && f[432] && !f[456] && f[436];
	assign leaf[12062] = !f[486] && f[432] && f[456] && !f[325];
	assign leaf[12063] = !f[486] && f[432] && f[456] && f[325];
	assign leaf[12064] = f[486] && !f[687] && !f[432] && !f[230];
	assign leaf[12065] = f[486] && !f[687] && !f[432] && f[230];
	assign leaf[12066] = f[486] && !f[687] && f[432] && !f[465];
	assign leaf[12067] = f[486] && !f[687] && f[432] && f[465];
	assign leaf[12068] = f[486] && f[687] && !f[548] && !f[690];
	assign leaf[12069] = f[486] && f[687] && !f[548] && f[690];
	assign leaf[12070] = f[486] && f[687] && f[548];
	
	// Tree 883, Classifier 3, Iteration: 88
	assign leaf[12071] = !f[429] && !f[491] && !f[461] && !f[407];
	assign leaf[12072] = !f[429] && !f[491] && !f[461] && f[407];
	assign leaf[12073] = !f[429] && !f[491] && f[461] && !f[544];
	assign leaf[12074] = !f[429] && !f[491] && f[461] && f[544];
	assign leaf[12075] = !f[429] && f[491] && !f[461] && !f[233];
	assign leaf[12076] = !f[429] && f[491] && !f[461] && f[233];
	assign leaf[12077] = !f[429] && f[491] && f[461] && !f[662];
	assign leaf[12078] = !f[429] && f[491] && f[461] && f[662];
	assign leaf[12079] = f[429] && !f[526] && !f[544] && !f[266];
	assign leaf[12080] = f[429] && !f[526] && !f[544] && f[266];
	assign leaf[12081] = f[429] && !f[526] && f[544] && !f[267];
	assign leaf[12082] = f[429] && !f[526] && f[544] && f[267];
	assign leaf[12083] = f[429] && f[526] && !f[521] && !f[317];
	assign leaf[12084] = f[429] && f[526] && !f[521] && f[317];
	assign leaf[12085] = f[429] && f[526] && f[521];
	
	// Tree 884, Classifier 4, Iteration: 88
	assign leaf[12086] = !f[465] && !f[424] && !f[380] && !f[439];
	assign leaf[12087] = !f[465] && !f[424] && !f[380] && f[439];
	assign leaf[12088] = !f[465] && !f[424] && f[380] && !f[466];
	assign leaf[12089] = !f[465] && !f[424] && f[380] && f[466];
	assign leaf[12090] = !f[465] && f[424];
	assign leaf[12091] = f[465] && !f[431] && !f[467] && !f[316];
	assign leaf[12092] = f[465] && !f[431] && !f[467] && f[316];
	assign leaf[12093] = f[465] && !f[431] && f[467] && !f[427];
	assign leaf[12094] = f[465] && !f[431] && f[467] && f[427];
	assign leaf[12095] = f[465] && f[431] && !f[216] && !f[286];
	assign leaf[12096] = f[465] && f[431] && !f[216] && f[286];
	assign leaf[12097] = f[465] && f[431] && f[216] && !f[184];
	assign leaf[12098] = f[465] && f[431] && f[216] && f[184];
	
	// Tree 885, Classifier 5, Iteration: 88
	assign leaf[12099] = !f[492] && !f[490] && !f[510] && !f[99];
	assign leaf[12100] = !f[492] && !f[490] && !f[510] && f[99];
	assign leaf[12101] = !f[492] && !f[490] && f[510] && !f[625];
	assign leaf[12102] = !f[492] && !f[490] && f[510] && f[625];
	assign leaf[12103] = !f[492] && f[490] && !f[261] && !f[331];
	assign leaf[12104] = !f[492] && f[490] && !f[261] && f[331];
	assign leaf[12105] = !f[492] && f[490] && f[261] && !f[319];
	assign leaf[12106] = !f[492] && f[490] && f[261] && f[319];
	assign leaf[12107] = f[492] && !f[625] && !f[511] && !f[684];
	assign leaf[12108] = f[492] && !f[625] && !f[511] && f[684];
	assign leaf[12109] = f[492] && !f[625] && f[511] && !f[538];
	assign leaf[12110] = f[492] && !f[625] && f[511] && f[538];
	assign leaf[12111] = f[492] && f[625] && !f[321] && !f[409];
	assign leaf[12112] = f[492] && f[625] && !f[321] && f[409];
	assign leaf[12113] = f[492] && f[625] && f[321] && !f[296];
	assign leaf[12114] = f[492] && f[625] && f[321] && f[296];
	
	// Tree 886, Classifier 6, Iteration: 88
	assign leaf[12115] = !f[629] && !f[383] && !f[549] && !f[521];
	assign leaf[12116] = !f[629] && !f[383] && !f[549] && f[521];
	assign leaf[12117] = !f[629] && !f[383] && f[549] && !f[514];
	assign leaf[12118] = !f[629] && !f[383] && f[549] && f[514];
	assign leaf[12119] = !f[629] && f[383] && !f[273] && !f[547];
	assign leaf[12120] = !f[629] && f[383] && !f[273] && f[547];
	assign leaf[12121] = !f[629] && f[383] && f[273];
	assign leaf[12122] = f[629] && !f[260] && !f[608] && !f[687];
	assign leaf[12123] = f[629] && !f[260] && !f[608] && f[687];
	assign leaf[12124] = f[629] && !f[260] && f[608] && !f[428];
	assign leaf[12125] = f[629] && !f[260] && f[608] && f[428];
	assign leaf[12126] = f[629] && f[260] && !f[464] && !f[545];
	assign leaf[12127] = f[629] && f[260] && !f[464] && f[545];
	assign leaf[12128] = f[629] && f[260] && f[464] && !f[483];
	assign leaf[12129] = f[629] && f[260] && f[464] && f[483];
	
	// Tree 887, Classifier 7, Iteration: 88
	assign leaf[12130] = !f[148] && !f[494] && !f[690] && !f[206];
	assign leaf[12131] = !f[148] && !f[494] && !f[690] && f[206];
	assign leaf[12132] = !f[148] && !f[494] && f[690] && !f[182];
	assign leaf[12133] = !f[148] && !f[494] && f[690] && f[182];
	assign leaf[12134] = !f[148] && f[494] && !f[346] && !f[185];
	assign leaf[12135] = !f[148] && f[494] && !f[346] && f[185];
	assign leaf[12136] = !f[148] && f[494] && f[346] && !f[407];
	assign leaf[12137] = !f[148] && f[494] && f[346] && f[407];
	assign leaf[12138] = f[148] && !f[356] && !f[211];
	assign leaf[12139] = f[148] && !f[356] && f[211] && !f[545];
	assign leaf[12140] = f[148] && !f[356] && f[211] && f[545];
	assign leaf[12141] = f[148] && f[356];
	
	// Tree 888, Classifier 8, Iteration: 88
	assign leaf[12142] = !f[678] && !f[161] && !f[570] && !f[632];
	assign leaf[12143] = !f[678] && !f[161] && !f[570] && f[632];
	assign leaf[12144] = !f[678] && !f[161] && f[570] && !f[572];
	assign leaf[12145] = !f[678] && !f[161] && f[570] && f[572];
	assign leaf[12146] = !f[678] && f[161] && !f[566] && !f[687];
	assign leaf[12147] = !f[678] && f[161] && !f[566] && f[687];
	assign leaf[12148] = !f[678] && f[161] && f[566] && !f[569];
	assign leaf[12149] = !f[678] && f[161] && f[566] && f[569];
	assign leaf[12150] = f[678] && !f[539] && !f[275];
	assign leaf[12151] = f[678] && !f[539] && f[275];
	assign leaf[12152] = f[678] && f[539];
	
	// Tree 889, Classifier 9, Iteration: 88
	assign leaf[12153] = !f[269] && !f[185] && !f[299] && !f[412];
	assign leaf[12154] = !f[269] && !f[185] && !f[299] && f[412];
	assign leaf[12155] = !f[269] && !f[185] && f[299] && !f[241];
	assign leaf[12156] = !f[269] && !f[185] && f[299] && f[241];
	assign leaf[12157] = !f[269] && f[185] && !f[212] && !f[657];
	assign leaf[12158] = !f[269] && f[185] && !f[212] && f[657];
	assign leaf[12159] = !f[269] && f[185] && f[212] && !f[156];
	assign leaf[12160] = !f[269] && f[185] && f[212] && f[156];
	assign leaf[12161] = f[269] && !f[187] && !f[322] && !f[486];
	assign leaf[12162] = f[269] && !f[187] && !f[322] && f[486];
	assign leaf[12163] = f[269] && !f[187] && f[322] && !f[403];
	assign leaf[12164] = f[269] && !f[187] && f[322] && f[403];
	assign leaf[12165] = f[269] && f[187] && !f[185] && !f[540];
	assign leaf[12166] = f[269] && f[187] && !f[185] && f[540];
	assign leaf[12167] = f[269] && f[187] && f[185] && !f[241];
	assign leaf[12168] = f[269] && f[187] && f[185] && f[241];
	
	// Tree 890, Classifier 0, Iteration: 89
	assign leaf[12169] = !f[602] && !f[456] && !f[687] && !f[356];
	assign leaf[12170] = !f[602] && !f[456] && !f[687] && f[356];
	assign leaf[12171] = !f[602] && !f[456] && f[687] && !f[156];
	assign leaf[12172] = !f[602] && !f[456] && f[687] && f[156];
	assign leaf[12173] = !f[602] && f[456] && !f[356] && !f[598];
	assign leaf[12174] = !f[602] && f[456] && !f[356] && f[598];
	assign leaf[12175] = !f[602] && f[456] && f[356] && !f[433];
	assign leaf[12176] = !f[602] && f[456] && f[356] && f[433];
	assign leaf[12177] = f[602] && !f[128] && !f[491] && !f[372];
	assign leaf[12178] = f[602] && !f[128] && !f[491] && f[372];
	assign leaf[12179] = f[602] && !f[128] && f[491] && !f[596];
	assign leaf[12180] = f[602] && !f[128] && f[491] && f[596];
	assign leaf[12181] = f[602] && f[128] && !f[322] && !f[435];
	assign leaf[12182] = f[602] && f[128] && !f[322] && f[435];
	assign leaf[12183] = f[602] && f[128] && f[322] && !f[463];
	assign leaf[12184] = f[602] && f[128] && f[322] && f[463];
	
	// Tree 891, Classifier 1, Iteration: 89
	assign leaf[12185] = !f[713] && !f[548] && !f[151] && !f[569];
	assign leaf[12186] = !f[713] && !f[548] && !f[151] && f[569];
	assign leaf[12187] = !f[713] && !f[548] && f[151] && !f[659];
	assign leaf[12188] = !f[713] && !f[548] && f[151] && f[659];
	assign leaf[12189] = !f[713] && f[548] && !f[576] && !f[129];
	assign leaf[12190] = !f[713] && f[548] && !f[576] && f[129];
	assign leaf[12191] = !f[713] && f[548] && f[576] && !f[405];
	assign leaf[12192] = !f[713] && f[548] && f[576] && f[405];
	assign leaf[12193] = f[713] && !f[349];
	assign leaf[12194] = f[713] && f[349];
	
	// Tree 892, Classifier 2, Iteration: 89
	assign leaf[12195] = !f[679] && !f[369] && !f[425] && !f[401];
	assign leaf[12196] = !f[679] && !f[369] && !f[425] && f[401];
	assign leaf[12197] = !f[679] && !f[369] && f[425] && !f[401];
	assign leaf[12198] = !f[679] && !f[369] && f[425] && f[401];
	assign leaf[12199] = !f[679] && f[369] && !f[490];
	assign leaf[12200] = !f[679] && f[369] && f[490] && !f[440];
	assign leaf[12201] = !f[679] && f[369] && f[490] && f[440];
	assign leaf[12202] = f[679] && !f[568] && !f[232];
	assign leaf[12203] = f[679] && !f[568] && f[232];
	assign leaf[12204] = f[679] && f[568] && !f[189];
	assign leaf[12205] = f[679] && f[568] && f[189];
	
	// Tree 893, Classifier 3, Iteration: 89
	assign leaf[12206] = !f[549] && !f[487] && !f[458] && !f[346];
	assign leaf[12207] = !f[549] && !f[487] && !f[458] && f[346];
	assign leaf[12208] = !f[549] && !f[487] && f[458] && !f[209];
	assign leaf[12209] = !f[549] && !f[487] && f[458] && f[209];
	assign leaf[12210] = !f[549] && f[487] && !f[457] && !f[511];
	assign leaf[12211] = !f[549] && f[487] && !f[457] && f[511];
	assign leaf[12212] = !f[549] && f[487] && f[457] && !f[206];
	assign leaf[12213] = !f[549] && f[487] && f[457] && f[206];
	assign leaf[12214] = f[549] && !f[657] && !f[439] && !f[542];
	assign leaf[12215] = f[549] && !f[657] && !f[439] && f[542];
	assign leaf[12216] = f[549] && !f[657] && f[439] && !f[493];
	assign leaf[12217] = f[549] && !f[657] && f[439] && f[493];
	assign leaf[12218] = f[549] && f[657] && !f[384] && !f[687];
	assign leaf[12219] = f[549] && f[657] && !f[384] && f[687];
	assign leaf[12220] = f[549] && f[657] && f[384] && !f[522];
	assign leaf[12221] = f[549] && f[657] && f[384] && f[522];
	
	// Tree 894, Classifier 4, Iteration: 89
	assign leaf[12222] = !f[303] && !f[386] && !f[234] && !f[684];
	assign leaf[12223] = !f[303] && !f[386] && !f[234] && f[684];
	assign leaf[12224] = !f[303] && !f[386] && f[234] && !f[237];
	assign leaf[12225] = !f[303] && !f[386] && f[234] && f[237];
	assign leaf[12226] = !f[303] && f[386] && !f[441] && !f[240];
	assign leaf[12227] = !f[303] && f[386] && !f[441] && f[240];
	assign leaf[12228] = !f[303] && f[386] && f[441] && !f[581];
	assign leaf[12229] = !f[303] && f[386] && f[441] && f[581];
	assign leaf[12230] = f[303] && !f[324] && !f[216] && !f[399];
	assign leaf[12231] = f[303] && !f[324] && !f[216] && f[399];
	assign leaf[12232] = f[303] && !f[324] && f[216];
	assign leaf[12233] = f[303] && f[324];
	
	// Tree 895, Classifier 5, Iteration: 89
	assign leaf[12234] = !f[351] && !f[454] && !f[296] && !f[327];
	assign leaf[12235] = !f[351] && !f[454] && !f[296] && f[327];
	assign leaf[12236] = !f[351] && !f[454] && f[296] && !f[184];
	assign leaf[12237] = !f[351] && !f[454] && f[296] && f[184];
	assign leaf[12238] = !f[351] && f[454] && !f[457] && !f[427];
	assign leaf[12239] = !f[351] && f[454] && !f[457] && f[427];
	assign leaf[12240] = !f[351] && f[454] && f[457] && !f[374];
	assign leaf[12241] = !f[351] && f[454] && f[457] && f[374];
	assign leaf[12242] = f[351] && !f[406] && !f[155] && !f[552];
	assign leaf[12243] = f[351] && !f[406] && !f[155] && f[552];
	assign leaf[12244] = f[351] && !f[406] && f[155] && !f[240];
	assign leaf[12245] = f[351] && !f[406] && f[155] && f[240];
	assign leaf[12246] = f[351] && f[406] && !f[540] && !f[348];
	assign leaf[12247] = f[351] && f[406] && !f[540] && f[348];
	assign leaf[12248] = f[351] && f[406] && f[540] && !f[325];
	assign leaf[12249] = f[351] && f[406] && f[540] && f[325];
	
	// Tree 896, Classifier 6, Iteration: 89
	assign leaf[12250] = !f[409] && !f[436] && !f[354] && !f[603];
	assign leaf[12251] = !f[409] && !f[436] && !f[354] && f[603];
	assign leaf[12252] = !f[409] && !f[436] && f[354] && !f[270];
	assign leaf[12253] = !f[409] && !f[436] && f[354] && f[270];
	assign leaf[12254] = !f[409] && f[436] && !f[576] && !f[440];
	assign leaf[12255] = !f[409] && f[436] && !f[576] && f[440];
	assign leaf[12256] = !f[409] && f[436] && f[576] && !f[406];
	assign leaf[12257] = !f[409] && f[436] && f[576] && f[406];
	assign leaf[12258] = f[409] && !f[435] && !f[326] && !f[429];
	assign leaf[12259] = f[409] && !f[435] && !f[326] && f[429];
	assign leaf[12260] = f[409] && !f[435] && f[326] && !f[239];
	assign leaf[12261] = f[409] && !f[435] && f[326] && f[239];
	assign leaf[12262] = f[409] && f[435] && !f[627] && !f[545];
	assign leaf[12263] = f[409] && f[435] && !f[627] && f[545];
	assign leaf[12264] = f[409] && f[435] && f[627] && !f[464];
	assign leaf[12265] = f[409] && f[435] && f[627] && f[464];
	
	// Tree 897, Classifier 7, Iteration: 89
	assign leaf[12266] = !f[510] && !f[428] && !f[457] && !f[544];
	assign leaf[12267] = !f[510] && !f[428] && !f[457] && f[544];
	assign leaf[12268] = !f[510] && !f[428] && f[457] && !f[401];
	assign leaf[12269] = !f[510] && !f[428] && f[457] && f[401];
	assign leaf[12270] = !f[510] && f[428] && !f[515] && !f[460];
	assign leaf[12271] = !f[510] && f[428] && !f[515] && f[460];
	assign leaf[12272] = !f[510] && f[428] && f[515] && !f[468];
	assign leaf[12273] = !f[510] && f[428] && f[515] && f[468];
	assign leaf[12274] = f[510] && !f[685] && !f[342];
	assign leaf[12275] = f[510] && !f[685] && f[342];
	assign leaf[12276] = f[510] && f[685];
	
	// Tree 898, Classifier 8, Iteration: 89
	assign leaf[12277] = !f[149] && !f[603] && !f[605] && !f[540];
	assign leaf[12278] = !f[149] && !f[603] && !f[605] && f[540];
	assign leaf[12279] = !f[149] && !f[603] && f[605] && !f[689];
	assign leaf[12280] = !f[149] && !f[603] && f[605] && f[689];
	assign leaf[12281] = !f[149] && f[603] && !f[604] && !f[630];
	assign leaf[12282] = !f[149] && f[603] && !f[604] && f[630];
	assign leaf[12283] = !f[149] && f[603] && f[604] && !f[427];
	assign leaf[12284] = !f[149] && f[603] && f[604] && f[427];
	assign leaf[12285] = f[149] && !f[204] && !f[465];
	assign leaf[12286] = f[149] && !f[204] && f[465] && !f[293];
	assign leaf[12287] = f[149] && !f[204] && f[465] && f[293];
	assign leaf[12288] = f[149] && f[204] && !f[319] && !f[239];
	assign leaf[12289] = f[149] && f[204] && !f[319] && f[239];
	assign leaf[12290] = f[149] && f[204] && f[319] && !f[344];
	assign leaf[12291] = f[149] && f[204] && f[319] && f[344];
	
	// Tree 899, Classifier 9, Iteration: 89
	assign leaf[12292] = !f[183] && !f[239] && !f[657] && !f[291];
	assign leaf[12293] = !f[183] && !f[239] && !f[657] && f[291];
	assign leaf[12294] = !f[183] && !f[239] && f[657] && !f[156];
	assign leaf[12295] = !f[183] && !f[239] && f[657] && f[156];
	assign leaf[12296] = !f[183] && f[239] && !f[433] && !f[381];
	assign leaf[12297] = !f[183] && f[239] && !f[433] && f[381];
	assign leaf[12298] = !f[183] && f[239] && f[433] && !f[462];
	assign leaf[12299] = !f[183] && f[239] && f[433] && f[462];
	assign leaf[12300] = f[183] && !f[211] && !f[398] && !f[184];
	assign leaf[12301] = f[183] && !f[211] && !f[398] && f[184];
	assign leaf[12302] = f[183] && !f[211] && f[398];
	assign leaf[12303] = f[183] && f[211] && !f[291] && !f[206];
	assign leaf[12304] = f[183] && f[211] && !f[291] && f[206];
	assign leaf[12305] = f[183] && f[211] && f[291] && !f[345];
	assign leaf[12306] = f[183] && f[211] && f[291] && f[345];
	
	// Tree 900, Classifier 0, Iteration: 90
	assign leaf[12307] = !f[240] && !f[325] && !f[214] && !f[331];
	assign leaf[12308] = !f[240] && !f[325] && !f[214] && f[331];
	assign leaf[12309] = !f[240] && !f[325] && f[214] && !f[128];
	assign leaf[12310] = !f[240] && !f[325] && f[214] && f[128];
	assign leaf[12311] = !f[240] && f[325] && !f[460] && !f[370];
	assign leaf[12312] = !f[240] && f[325] && !f[460] && f[370];
	assign leaf[12313] = !f[240] && f[325] && f[460];
	assign leaf[12314] = f[240] && !f[466] && !f[374] && !f[511];
	assign leaf[12315] = f[240] && !f[466] && !f[374] && f[511];
	assign leaf[12316] = f[240] && !f[466] && f[374] && !f[468];
	assign leaf[12317] = f[240] && !f[466] && f[374] && f[468];
	assign leaf[12318] = f[240] && f[466] && !f[403] && !f[400];
	assign leaf[12319] = f[240] && f[466] && !f[403] && f[400];
	assign leaf[12320] = f[240] && f[466] && f[403] && !f[457];
	assign leaf[12321] = f[240] && f[466] && f[403] && f[457];
	
	// Tree 901, Classifier 1, Iteration: 90
	assign leaf[12322] = !f[712] && !f[440] && !f[578] && !f[177];
	assign leaf[12323] = !f[712] && !f[440] && !f[578] && f[177];
	assign leaf[12324] = !f[712] && !f[440] && f[578] && !f[517];
	assign leaf[12325] = !f[712] && !f[440] && f[578] && f[517];
	assign leaf[12326] = !f[712] && f[440];
	assign leaf[12327] = f[712] && !f[432];
	assign leaf[12328] = f[712] && f[432];
	
	// Tree 902, Classifier 2, Iteration: 90
	assign leaf[12329] = !f[570] && !f[480] && !f[268] && !f[180];
	assign leaf[12330] = !f[570] && !f[480] && !f[268] && f[180];
	assign leaf[12331] = !f[570] && !f[480] && f[268] && !f[458];
	assign leaf[12332] = !f[570] && !f[480] && f[268] && f[458];
	assign leaf[12333] = !f[570] && f[480] && !f[461];
	assign leaf[12334] = !f[570] && f[480] && f[461];
	assign leaf[12335] = f[570] && !f[655] && !f[489] && !f[458];
	assign leaf[12336] = f[570] && !f[655] && !f[489] && f[458];
	assign leaf[12337] = f[570] && !f[655] && f[489] && !f[681];
	assign leaf[12338] = f[570] && !f[655] && f[489] && f[681];
	assign leaf[12339] = f[570] && f[655] && !f[403] && !f[406];
	assign leaf[12340] = f[570] && f[655] && !f[403] && f[406];
	assign leaf[12341] = f[570] && f[655] && f[403] && !f[484];
	assign leaf[12342] = f[570] && f[655] && f[403] && f[484];
	
	// Tree 903, Classifier 3, Iteration: 90
	assign leaf[12343] = !f[492] && !f[547] && !f[517] && !f[322];
	assign leaf[12344] = !f[492] && !f[547] && !f[517] && f[322];
	assign leaf[12345] = !f[492] && !f[547] && f[517] && !f[572];
	assign leaf[12346] = !f[492] && !f[547] && f[517] && f[572];
	assign leaf[12347] = !f[492] && f[547] && !f[554] && !f[381];
	assign leaf[12348] = !f[492] && f[547] && !f[554] && f[381];
	assign leaf[12349] = !f[492] && f[547] && f[554] && !f[436];
	assign leaf[12350] = !f[492] && f[547] && f[554] && f[436];
	assign leaf[12351] = f[492] && !f[437] && !f[354] && !f[404];
	assign leaf[12352] = f[492] && !f[437] && !f[354] && f[404];
	assign leaf[12353] = f[492] && !f[437] && f[354] && !f[483];
	assign leaf[12354] = f[492] && !f[437] && f[354] && f[483];
	assign leaf[12355] = f[492] && f[437] && !f[625] && !f[274];
	assign leaf[12356] = f[492] && f[437] && !f[625] && f[274];
	assign leaf[12357] = f[492] && f[437] && f[625] && !f[154];
	assign leaf[12358] = f[492] && f[437] && f[625] && f[154];
	
	// Tree 904, Classifier 4, Iteration: 90
	assign leaf[12359] = !f[389] && !f[128] && !f[555] && !f[370];
	assign leaf[12360] = !f[389] && !f[128] && !f[555] && f[370];
	assign leaf[12361] = !f[389] && !f[128] && f[555] && !f[466];
	assign leaf[12362] = !f[389] && !f[128] && f[555] && f[466];
	assign leaf[12363] = !f[389] && f[128] && !f[497] && !f[376];
	assign leaf[12364] = !f[389] && f[128] && !f[497] && f[376];
	assign leaf[12365] = !f[389] && f[128] && f[497] && !f[293];
	assign leaf[12366] = !f[389] && f[128] && f[497] && f[293];
	assign leaf[12367] = f[389];
	
	// Tree 905, Classifier 5, Iteration: 90
	assign leaf[12368] = !f[119] && !f[322] && !f[519] && !f[517];
	assign leaf[12369] = !f[119] && !f[322] && !f[519] && f[517];
	assign leaf[12370] = !f[119] && !f[322] && f[519] && !f[295];
	assign leaf[12371] = !f[119] && !f[322] && f[519] && f[295];
	assign leaf[12372] = !f[119] && f[322] && !f[491] && !f[462];
	assign leaf[12373] = !f[119] && f[322] && !f[491] && f[462];
	assign leaf[12374] = !f[119] && f[322] && f[491] && !f[265];
	assign leaf[12375] = !f[119] && f[322] && f[491] && f[265];
	assign leaf[12376] = f[119] && !f[609];
	assign leaf[12377] = f[119] && f[609];
	
	// Tree 906, Classifier 6, Iteration: 90
	assign leaf[12378] = !f[355] && !f[272] && !f[297] && !f[358];
	assign leaf[12379] = !f[355] && !f[272] && !f[297] && f[358];
	assign leaf[12380] = !f[355] && !f[272] && f[297] && !f[625];
	assign leaf[12381] = !f[355] && !f[272] && f[297] && f[625];
	assign leaf[12382] = !f[355] && f[272] && !f[635] && !f[291];
	assign leaf[12383] = !f[355] && f[272] && !f[635] && f[291];
	assign leaf[12384] = !f[355] && f[272] && f[635];
	assign leaf[12385] = f[355] && !f[352] && !f[441] && !f[358];
	assign leaf[12386] = f[355] && !f[352] && !f[441] && f[358];
	assign leaf[12387] = f[355] && !f[352] && f[441] && !f[456];
	assign leaf[12388] = f[355] && !f[352] && f[441] && f[456];
	assign leaf[12389] = f[355] && f[352] && !f[349] && !f[239];
	assign leaf[12390] = f[355] && f[352] && !f[349] && f[239];
	assign leaf[12391] = f[355] && f[352] && f[349] && !f[400];
	assign leaf[12392] = f[355] && f[352] && f[349] && f[400];
	
	// Tree 907, Classifier 7, Iteration: 90
	assign leaf[12393] = !f[704] && !f[595] && !f[720] && !f[206];
	assign leaf[12394] = !f[704] && !f[595] && !f[720] && f[206];
	assign leaf[12395] = !f[704] && !f[595] && f[720] && !f[266];
	assign leaf[12396] = !f[704] && !f[595] && f[720] && f[266];
	assign leaf[12397] = !f[704] && f[595] && !f[573] && !f[434];
	assign leaf[12398] = !f[704] && f[595] && !f[573] && f[434];
	assign leaf[12399] = !f[704] && f[595] && f[573] && !f[294];
	assign leaf[12400] = !f[704] && f[595] && f[573] && f[294];
	assign leaf[12401] = f[704];
	
	// Tree 908, Classifier 8, Iteration: 90
	assign leaf[12402] = !f[486] && !f[488] && !f[517] && !f[456];
	assign leaf[12403] = !f[486] && !f[488] && !f[517] && f[456];
	assign leaf[12404] = !f[486] && !f[488] && f[517] && !f[549];
	assign leaf[12405] = !f[486] && !f[488] && f[517] && f[549];
	assign leaf[12406] = !f[486] && f[488] && !f[352] && !f[489];
	assign leaf[12407] = !f[486] && f[488] && !f[352] && f[489];
	assign leaf[12408] = !f[486] && f[488] && f[352] && !f[290];
	assign leaf[12409] = !f[486] && f[488] && f[352] && f[290];
	assign leaf[12410] = f[486] && !f[516] && !f[541] && !f[543];
	assign leaf[12411] = f[486] && !f[516] && !f[541] && f[543];
	assign leaf[12412] = f[486] && !f[516] && f[541] && !f[462];
	assign leaf[12413] = f[486] && !f[516] && f[541] && f[462];
	assign leaf[12414] = f[486] && f[516] && !f[400] && !f[512];
	assign leaf[12415] = f[486] && f[516] && !f[400] && f[512];
	assign leaf[12416] = f[486] && f[516] && f[400] && !f[513];
	assign leaf[12417] = f[486] && f[516] && f[400] && f[513];
	
	// Tree 909, Classifier 9, Iteration: 90
	assign leaf[12418] = !f[256] && !f[342] && !f[387] && !f[320];
	assign leaf[12419] = !f[256] && !f[342] && !f[387] && f[320];
	assign leaf[12420] = !f[256] && !f[342] && f[387];
	assign leaf[12421] = !f[256] && f[342] && !f[290] && !f[687];
	assign leaf[12422] = !f[256] && f[342] && !f[290] && f[687];
	assign leaf[12423] = !f[256] && f[342] && f[290] && !f[454];
	assign leaf[12424] = !f[256] && f[342] && f[290] && f[454];
	assign leaf[12425] = f[256] && !f[398];
	assign leaf[12426] = f[256] && f[398];
	
	// Tree 910, Classifier 0, Iteration: 91
	assign leaf[12427] = !f[663] && !f[583] && !f[513] && !f[328];
	assign leaf[12428] = !f[663] && !f[583] && !f[513] && f[328];
	assign leaf[12429] = !f[663] && !f[583] && f[513] && !f[183];
	assign leaf[12430] = !f[663] && !f[583] && f[513] && f[183];
	assign leaf[12431] = !f[663] && f[583];
	assign leaf[12432] = f[663] && !f[346];
	assign leaf[12433] = f[663] && f[346];
	
	// Tree 911, Classifier 1, Iteration: 91
	assign leaf[12434] = !f[215] && !f[381] && !f[241] && !f[210];
	assign leaf[12435] = !f[215] && !f[381] && !f[241] && f[210];
	assign leaf[12436] = !f[215] && !f[381] && f[241] && !f[575];
	assign leaf[12437] = !f[215] && !f[381] && f[241] && f[575];
	assign leaf[12438] = !f[215] && f[381] && !f[548] && !f[240];
	assign leaf[12439] = !f[215] && f[381] && !f[548] && f[240];
	assign leaf[12440] = !f[215] && f[381] && f[548] && !f[346];
	assign leaf[12441] = !f[215] && f[381] && f[548] && f[346];
	assign leaf[12442] = f[215] && !f[324];
	assign leaf[12443] = f[215] && f[324] && !f[381] && !f[519];
	assign leaf[12444] = f[215] && f[324] && !f[381] && f[519];
	assign leaf[12445] = f[215] && f[324] && f[381] && !f[209];
	assign leaf[12446] = f[215] && f[324] && f[381] && f[209];
	
	// Tree 912, Classifier 2, Iteration: 91
	assign leaf[12447] = !f[512] && !f[575] && !f[714] && !f[654];
	assign leaf[12448] = !f[512] && !f[575] && !f[714] && f[654];
	assign leaf[12449] = !f[512] && !f[575] && f[714];
	assign leaf[12450] = !f[512] && f[575] && !f[403] && !f[100];
	assign leaf[12451] = !f[512] && f[575] && !f[403] && f[100];
	assign leaf[12452] = !f[512] && f[575] && f[403] && !f[427];
	assign leaf[12453] = !f[512] && f[575] && f[403] && f[427];
	assign leaf[12454] = f[512] && !f[433] && !f[233] && !f[265];
	assign leaf[12455] = f[512] && !f[433] && !f[233] && f[265];
	assign leaf[12456] = f[512] && !f[433] && f[233] && !f[595];
	assign leaf[12457] = f[512] && !f[433] && f[233] && f[595];
	assign leaf[12458] = f[512] && f[433] && !f[457] && !f[186];
	assign leaf[12459] = f[512] && f[433] && !f[457] && f[186];
	assign leaf[12460] = f[512] && f[433] && f[457] && !f[245];
	assign leaf[12461] = f[512] && f[433] && f[457] && f[245];
	
	// Tree 913, Classifier 3, Iteration: 91
	assign leaf[12462] = !f[427] && !f[705] && !f[591] && !f[218];
	assign leaf[12463] = !f[427] && !f[705] && !f[591] && f[218];
	assign leaf[12464] = !f[427] && !f[705] && f[591] && !f[159];
	assign leaf[12465] = !f[427] && !f[705] && f[591] && f[159];
	assign leaf[12466] = !f[427] && f[705];
	assign leaf[12467] = f[427] && !f[219] && !f[212] && !f[204];
	assign leaf[12468] = f[427] && !f[219] && !f[212] && f[204];
	assign leaf[12469] = f[427] && !f[219] && f[212] && !f[429];
	assign leaf[12470] = f[427] && !f[219] && f[212] && f[429];
	assign leaf[12471] = f[427] && f[219];
	
	// Tree 914, Classifier 4, Iteration: 91
	assign leaf[12472] = !f[746] && !f[400] && !f[490] && !f[628];
	assign leaf[12473] = !f[746] && !f[400] && !f[490] && f[628];
	assign leaf[12474] = !f[746] && !f[400] && f[490] && !f[376];
	assign leaf[12475] = !f[746] && !f[400] && f[490] && f[376];
	assign leaf[12476] = !f[746] && f[400] && !f[547] && !f[658];
	assign leaf[12477] = !f[746] && f[400] && !f[547] && f[658];
	assign leaf[12478] = !f[746] && f[400] && f[547] && !f[549];
	assign leaf[12479] = !f[746] && f[400] && f[547] && f[549];
	assign leaf[12480] = f[746];
	
	// Tree 915, Classifier 5, Iteration: 91
	assign leaf[12481] = !f[485] && !f[291] && !f[596] && !f[266];
	assign leaf[12482] = !f[485] && !f[291] && !f[596] && f[266];
	assign leaf[12483] = !f[485] && !f[291] && f[596] && !f[235];
	assign leaf[12484] = !f[485] && !f[291] && f[596] && f[235];
	assign leaf[12485] = !f[485] && f[291] && !f[207] && !f[407];
	assign leaf[12486] = !f[485] && f[291] && !f[207] && f[407];
	assign leaf[12487] = !f[485] && f[291] && f[207] && !f[235];
	assign leaf[12488] = !f[485] && f[291] && f[207] && f[235];
	assign leaf[12489] = f[485] && !f[407] && !f[136] && !f[541];
	assign leaf[12490] = f[485] && !f[407] && !f[136] && f[541];
	assign leaf[12491] = f[485] && !f[407] && f[136];
	assign leaf[12492] = f[485] && f[407] && !f[515] && !f[569];
	assign leaf[12493] = f[485] && f[407] && !f[515] && f[569];
	assign leaf[12494] = f[485] && f[407] && f[515] && !f[577];
	assign leaf[12495] = f[485] && f[407] && f[515] && f[577];
	
	// Tree 916, Classifier 6, Iteration: 91
	assign leaf[12496] = !f[516] && !f[485] && !f[483] && !f[486];
	assign leaf[12497] = !f[516] && !f[485] && !f[483] && f[486];
	assign leaf[12498] = !f[516] && !f[485] && f[483] && !f[497];
	assign leaf[12499] = !f[516] && !f[485] && f[483] && f[497];
	assign leaf[12500] = !f[516] && f[485] && !f[373] && !f[262];
	assign leaf[12501] = !f[516] && f[485] && !f[373] && f[262];
	assign leaf[12502] = !f[516] && f[485] && f[373] && !f[241];
	assign leaf[12503] = !f[516] && f[485] && f[373] && f[241];
	assign leaf[12504] = f[516] && !f[275] && !f[216] && !f[294];
	assign leaf[12505] = f[516] && !f[275] && !f[216] && f[294];
	assign leaf[12506] = f[516] && !f[275] && f[216] && !f[380];
	assign leaf[12507] = f[516] && !f[275] && f[216] && f[380];
	assign leaf[12508] = f[516] && f[275];
	
	// Tree 917, Classifier 7, Iteration: 91
	assign leaf[12509] = !f[148] && !f[312] && !f[463] && !f[601];
	assign leaf[12510] = !f[148] && !f[312] && !f[463] && f[601];
	assign leaf[12511] = !f[148] && !f[312] && f[463] && !f[578];
	assign leaf[12512] = !f[148] && !f[312] && f[463] && f[578];
	assign leaf[12513] = !f[148] && f[312] && !f[553] && !f[398];
	assign leaf[12514] = !f[148] && f[312] && !f[553] && f[398];
	assign leaf[12515] = !f[148] && f[312] && f[553];
	assign leaf[12516] = f[148] && !f[630] && !f[184];
	assign leaf[12517] = f[148] && !f[630] && f[184];
	assign leaf[12518] = f[148] && f[630] && !f[655];
	assign leaf[12519] = f[148] && f[630] && f[655];
	
	// Tree 918, Classifier 8, Iteration: 91
	assign leaf[12520] = !f[440] && !f[388] && !f[315] && !f[410];
	assign leaf[12521] = !f[440] && !f[388] && !f[315] && f[410];
	assign leaf[12522] = !f[440] && !f[388] && f[315] && !f[292];
	assign leaf[12523] = !f[440] && !f[388] && f[315] && f[292];
	assign leaf[12524] = !f[440] && f[388];
	assign leaf[12525] = f[440] && !f[555] && !f[625] && !f[381];
	assign leaf[12526] = f[440] && !f[555] && !f[625] && f[381];
	assign leaf[12527] = f[440] && !f[555] && f[625] && !f[458];
	assign leaf[12528] = f[440] && !f[555] && f[625] && f[458];
	assign leaf[12529] = f[440] && f[555] && !f[525];
	assign leaf[12530] = f[440] && f[555] && f[525] && !f[354];
	assign leaf[12531] = f[440] && f[555] && f[525] && f[354];
	
	// Tree 919, Classifier 9, Iteration: 91
	assign leaf[12532] = !f[742] && !f[740] && !f[182] && !f[266];
	assign leaf[12533] = !f[742] && !f[740] && !f[182] && f[266];
	assign leaf[12534] = !f[742] && !f[740] && f[182] && !f[237];
	assign leaf[12535] = !f[742] && !f[740] && f[182] && f[237];
	assign leaf[12536] = !f[742] && f[740] && !f[406] && !f[461];
	assign leaf[12537] = !f[742] && f[740] && !f[406] && f[461];
	assign leaf[12538] = !f[742] && f[740] && f[406] && !f[289];
	assign leaf[12539] = !f[742] && f[740] && f[406] && f[289];
	assign leaf[12540] = f[742] && !f[326] && !f[319];
	assign leaf[12541] = f[742] && !f[326] && f[319];
	assign leaf[12542] = f[742] && f[326] && !f[601] && !f[458];
	assign leaf[12543] = f[742] && f[326] && !f[601] && f[458];
	assign leaf[12544] = f[742] && f[326] && f[601];
	
	// Tree 920, Classifier 0, Iteration: 92
	assign leaf[12545] = !f[605] && !f[260] && !f[242] && !f[566];
	assign leaf[12546] = !f[605] && !f[260] && !f[242] && f[566];
	assign leaf[12547] = !f[605] && !f[260] && f[242] && !f[683];
	assign leaf[12548] = !f[605] && !f[260] && f[242] && f[683];
	assign leaf[12549] = !f[605] && f[260] && !f[359] && !f[545];
	assign leaf[12550] = !f[605] && f[260] && !f[359] && f[545];
	assign leaf[12551] = !f[605] && f[260] && f[359];
	assign leaf[12552] = f[605] && !f[397] && !f[597] && !f[599];
	assign leaf[12553] = f[605] && !f[397] && !f[597] && f[599];
	assign leaf[12554] = f[605] && !f[397] && f[597] && !f[484];
	assign leaf[12555] = f[605] && !f[397] && f[597] && f[484];
	assign leaf[12556] = f[605] && f[397] && !f[207];
	assign leaf[12557] = f[605] && f[397] && f[207] && !f[428];
	assign leaf[12558] = f[605] && f[397] && f[207] && f[428];
	
	// Tree 921, Classifier 1, Iteration: 92
	assign leaf[12559] = !f[95] && !f[609] && !f[708] && !f[204];
	assign leaf[12560] = !f[95] && !f[609] && !f[708] && f[204];
	assign leaf[12561] = !f[95] && !f[609] && f[708];
	assign leaf[12562] = !f[95] && f[609] && !f[516];
	assign leaf[12563] = !f[95] && f[609] && f[516];
	assign leaf[12564] = f[95];
	
	// Tree 922, Classifier 2, Iteration: 92
	assign leaf[12565] = !f[455] && !f[611] && !f[430] && !f[346];
	assign leaf[12566] = !f[455] && !f[611] && !f[430] && f[346];
	assign leaf[12567] = !f[455] && !f[611] && f[430] && !f[484];
	assign leaf[12568] = !f[455] && !f[611] && f[430] && f[484];
	assign leaf[12569] = !f[455] && f[611] && !f[210];
	assign leaf[12570] = !f[455] && f[611] && f[210];
	assign leaf[12571] = f[455] && !f[261] && !f[573] && !f[406];
	assign leaf[12572] = f[455] && !f[261] && !f[573] && f[406];
	assign leaf[12573] = f[455] && !f[261] && f[573] && !f[154];
	assign leaf[12574] = f[455] && !f[261] && f[573] && f[154];
	assign leaf[12575] = f[455] && f[261] && !f[566] && !f[402];
	assign leaf[12576] = f[455] && f[261] && !f[566] && f[402];
	assign leaf[12577] = f[455] && f[261] && f[566] && !f[158];
	assign leaf[12578] = f[455] && f[261] && f[566] && f[158];
	
	// Tree 923, Classifier 3, Iteration: 92
	assign leaf[12579] = !f[637] && !f[555] && !f[122] && !f[347];
	assign leaf[12580] = !f[637] && !f[555] && !f[122] && f[347];
	assign leaf[12581] = !f[637] && !f[555] && f[122] && !f[233];
	assign leaf[12582] = !f[637] && !f[555] && f[122] && f[233];
	assign leaf[12583] = !f[637] && f[555] && !f[320];
	assign leaf[12584] = !f[637] && f[555] && f[320] && !f[597];
	assign leaf[12585] = !f[637] && f[555] && f[320] && f[597];
	assign leaf[12586] = f[637] && !f[207] && !f[211];
	assign leaf[12587] = f[637] && !f[207] && f[211];
	assign leaf[12588] = f[637] && f[207] && !f[607] && !f[177];
	assign leaf[12589] = f[637] && f[207] && !f[607] && f[177];
	assign leaf[12590] = f[637] && f[207] && f[607] && !f[321];
	assign leaf[12591] = f[637] && f[207] && f[607] && f[321];
	
	// Tree 924, Classifier 4, Iteration: 92
	assign leaf[12592] = !f[494] && !f[435] && !f[520] && !f[408];
	assign leaf[12593] = !f[494] && !f[435] && !f[520] && f[408];
	assign leaf[12594] = !f[494] && !f[435] && f[520] && !f[295];
	assign leaf[12595] = !f[494] && !f[435] && f[520] && f[295];
	assign leaf[12596] = !f[494] && f[435] && !f[238] && !f[264];
	assign leaf[12597] = !f[494] && f[435] && !f[238] && f[264];
	assign leaf[12598] = !f[494] && f[435] && f[238] && !f[294];
	assign leaf[12599] = !f[494] && f[435] && f[238] && f[294];
	assign leaf[12600] = f[494] && !f[434] && !f[350] && !f[600];
	assign leaf[12601] = f[494] && !f[434] && !f[350] && f[600];
	assign leaf[12602] = f[494] && !f[434] && f[350] && !f[635];
	assign leaf[12603] = f[494] && !f[434] && f[350] && f[635];
	assign leaf[12604] = f[494] && f[434] && !f[510] && !f[454];
	assign leaf[12605] = f[494] && f[434] && !f[510] && f[454];
	assign leaf[12606] = f[494] && f[434] && f[510] && !f[498];
	assign leaf[12607] = f[494] && f[434] && f[510] && f[498];
	
	// Tree 925, Classifier 5, Iteration: 92
	assign leaf[12608] = !f[627] && !f[428] && !f[271] && !f[184];
	assign leaf[12609] = !f[627] && !f[428] && !f[271] && f[184];
	assign leaf[12610] = !f[627] && !f[428] && f[271] && !f[269];
	assign leaf[12611] = !f[627] && !f[428] && f[271] && f[269];
	assign leaf[12612] = !f[627] && f[428] && !f[290] && !f[510];
	assign leaf[12613] = !f[627] && f[428] && !f[290] && f[510];
	assign leaf[12614] = !f[627] && f[428] && f[290] && !f[128];
	assign leaf[12615] = !f[627] && f[428] && f[290] && f[128];
	assign leaf[12616] = f[627] && !f[463] && !f[234] && !f[290];
	assign leaf[12617] = f[627] && !f[463] && !f[234] && f[290];
	assign leaf[12618] = f[627] && !f[463] && f[234] && !f[269];
	assign leaf[12619] = f[627] && !f[463] && f[234] && f[269];
	assign leaf[12620] = f[627] && f[463] && !f[547] && !f[321];
	assign leaf[12621] = f[627] && f[463] && !f[547] && f[321];
	assign leaf[12622] = f[627] && f[463] && f[547] && !f[384];
	assign leaf[12623] = f[627] && f[463] && f[547] && f[384];
	
	// Tree 926, Classifier 6, Iteration: 92
	assign leaf[12624] = !f[522] && !f[570] && !f[634] && !f[242];
	assign leaf[12625] = !f[522] && !f[570] && !f[634] && f[242];
	assign leaf[12626] = !f[522] && !f[570] && f[634] && !f[184];
	assign leaf[12627] = !f[522] && !f[570] && f[634] && f[184];
	assign leaf[12628] = !f[522] && f[570] && !f[408] && !f[434];
	assign leaf[12629] = !f[522] && f[570] && !f[408] && f[434];
	assign leaf[12630] = !f[522] && f[570] && f[408] && !f[466];
	assign leaf[12631] = !f[522] && f[570] && f[408] && f[466];
	assign leaf[12632] = f[522] && !f[261] && !f[151] && !f[217];
	assign leaf[12633] = f[522] && !f[261] && !f[151] && f[217];
	assign leaf[12634] = f[522] && !f[261] && f[151] && !f[239];
	assign leaf[12635] = f[522] && !f[261] && f[151] && f[239];
	assign leaf[12636] = f[522] && f[261] && !f[264] && !f[459];
	assign leaf[12637] = f[522] && f[261] && !f[264] && f[459];
	assign leaf[12638] = f[522] && f[261] && f[264] && !f[125];
	assign leaf[12639] = f[522] && f[261] && f[264] && f[125];
	
	// Tree 927, Classifier 7, Iteration: 92
	assign leaf[12640] = !f[298] && !f[323] && !f[287] && !f[715];
	assign leaf[12641] = !f[298] && !f[323] && !f[287] && f[715];
	assign leaf[12642] = !f[298] && !f[323] && f[287] && !f[461];
	assign leaf[12643] = !f[298] && !f[323] && f[287] && f[461];
	assign leaf[12644] = !f[298] && f[323] && !f[687] && !f[431];
	assign leaf[12645] = !f[298] && f[323] && !f[687] && f[431];
	assign leaf[12646] = !f[298] && f[323] && f[687] && !f[347];
	assign leaf[12647] = !f[298] && f[323] && f[687] && f[347];
	assign leaf[12648] = f[298] && !f[406] && !f[158] && !f[351];
	assign leaf[12649] = f[298] && !f[406] && !f[158] && f[351];
	assign leaf[12650] = f[298] && !f[406] && f[158];
	assign leaf[12651] = f[298] && f[406] && !f[570] && !f[202];
	assign leaf[12652] = f[298] && f[406] && !f[570] && f[202];
	assign leaf[12653] = f[298] && f[406] && f[570] && !f[602];
	assign leaf[12654] = f[298] && f[406] && f[570] && f[602];
	
	// Tree 928, Classifier 8, Iteration: 92
	assign leaf[12655] = !f[275] && !f[679] && !f[457] && !f[597];
	assign leaf[12656] = !f[275] && !f[679] && !f[457] && f[597];
	assign leaf[12657] = !f[275] && !f[679] && f[457] && !f[488];
	assign leaf[12658] = !f[275] && !f[679] && f[457] && f[488];
	assign leaf[12659] = !f[275] && f[679] && !f[540] && !f[378];
	assign leaf[12660] = !f[275] && f[679] && !f[540] && f[378];
	assign leaf[12661] = !f[275] && f[679] && f[540] && !f[625];
	assign leaf[12662] = !f[275] && f[679] && f[540] && f[625];
	assign leaf[12663] = f[275] && !f[520] && !f[457] && !f[214];
	assign leaf[12664] = f[275] && !f[520] && !f[457] && f[214];
	assign leaf[12665] = f[275] && !f[520] && f[457] && !f[485];
	assign leaf[12666] = f[275] && !f[520] && f[457] && f[485];
	assign leaf[12667] = f[275] && f[520] && !f[207] && !f[466];
	assign leaf[12668] = f[275] && f[520] && !f[207] && f[466];
	assign leaf[12669] = f[275] && f[520] && f[207] && !f[514];
	assign leaf[12670] = f[275] && f[520] && f[207] && f[514];
	
	// Tree 929, Classifier 9, Iteration: 92
	assign leaf[12671] = !f[740] && !f[472] && !f[184] && !f[602];
	assign leaf[12672] = !f[740] && !f[472] && !f[184] && f[602];
	assign leaf[12673] = !f[740] && !f[472] && f[184] && !f[717];
	assign leaf[12674] = !f[740] && !f[472] && f[184] && f[717];
	assign leaf[12675] = !f[740] && f[472];
	assign leaf[12676] = f[740] && !f[544] && !f[490] && !f[290];
	assign leaf[12677] = f[740] && !f[544] && !f[490] && f[290];
	assign leaf[12678] = f[740] && !f[544] && f[490] && !f[713];
	assign leaf[12679] = f[740] && !f[544] && f[490] && f[713];
	assign leaf[12680] = f[740] && f[544];
	
	// Tree 930, Classifier 0, Iteration: 93
	assign leaf[12681] = !f[294] && !f[351] && !f[518] && !f[344];
	assign leaf[12682] = !f[294] && !f[351] && !f[518] && f[344];
	assign leaf[12683] = !f[294] && !f[351] && f[518] && !f[455];
	assign leaf[12684] = !f[294] && !f[351] && f[518] && f[455];
	assign leaf[12685] = !f[294] && f[351] && !f[376];
	assign leaf[12686] = !f[294] && f[351] && f[376];
	assign leaf[12687] = f[294] && !f[99] && !f[384] && !f[160];
	assign leaf[12688] = f[294] && !f[99] && !f[384] && f[160];
	assign leaf[12689] = f[294] && !f[99] && f[384] && !f[402];
	assign leaf[12690] = f[294] && !f[99] && f[384] && f[402];
	assign leaf[12691] = f[294] && f[99];
	
	// Tree 931, Classifier 1, Iteration: 93
	assign leaf[12692] = !f[715] && !f[712] && !f[374] && !f[244];
	assign leaf[12693] = !f[715] && !f[712] && !f[374] && f[244];
	assign leaf[12694] = !f[715] && !f[712] && f[374] && !f[323];
	assign leaf[12695] = !f[715] && !f[712] && f[374] && f[323];
	assign leaf[12696] = !f[715] && f[712] && !f[376];
	assign leaf[12697] = !f[715] && f[712] && f[376];
	assign leaf[12698] = f[715] && !f[346];
	assign leaf[12699] = f[715] && f[346];
	
	// Tree 932, Classifier 2, Iteration: 93
	assign leaf[12700] = !f[598] && !f[655] && !f[208] && !f[635];
	assign leaf[12701] = !f[598] && !f[655] && !f[208] && f[635];
	assign leaf[12702] = !f[598] && !f[655] && f[208] && !f[238];
	assign leaf[12703] = !f[598] && !f[655] && f[208] && f[238];
	assign leaf[12704] = !f[598] && f[655] && !f[688] && !f[607];
	assign leaf[12705] = !f[598] && f[655] && !f[688] && f[607];
	assign leaf[12706] = !f[598] && f[655] && f[688];
	assign leaf[12707] = f[598] && !f[179] && !f[272] && !f[97];
	assign leaf[12708] = f[598] && !f[179] && !f[272] && f[97];
	assign leaf[12709] = f[598] && !f[179] && f[272] && !f[264];
	assign leaf[12710] = f[598] && !f[179] && f[272] && f[264];
	assign leaf[12711] = f[598] && f[179] && !f[268] && !f[409];
	assign leaf[12712] = f[598] && f[179] && !f[268] && f[409];
	assign leaf[12713] = f[598] && f[179] && f[268] && !f[432];
	assign leaf[12714] = f[598] && f[179] && f[268] && f[432];
	
	// Tree 933, Classifier 3, Iteration: 93
	assign leaf[12715] = !f[342] && !f[260] && !f[177] && !f[574];
	assign leaf[12716] = !f[342] && !f[260] && !f[177] && f[574];
	assign leaf[12717] = !f[342] && !f[260] && f[177] && !f[347];
	assign leaf[12718] = !f[342] && !f[260] && f[177] && f[347];
	assign leaf[12719] = !f[342] && f[260] && !f[289] && !f[347];
	assign leaf[12720] = !f[342] && f[260] && !f[289] && f[347];
	assign leaf[12721] = !f[342] && f[260] && f[289] && !f[236];
	assign leaf[12722] = !f[342] && f[260] && f[289] && f[236];
	assign leaf[12723] = f[342] && !f[323] && !f[355];
	assign leaf[12724] = f[342] && !f[323] && f[355] && !f[634];
	assign leaf[12725] = f[342] && !f[323] && f[355] && f[634];
	assign leaf[12726] = f[342] && f[323] && !f[525];
	assign leaf[12727] = f[342] && f[323] && f[525] && !f[270];
	assign leaf[12728] = f[342] && f[323] && f[525] && f[270];
	
	// Tree 934, Classifier 4, Iteration: 93
	assign leaf[12729] = !f[237] && !f[261] && !f[239] && !f[236];
	assign leaf[12730] = !f[237] && !f[261] && !f[239] && f[236];
	assign leaf[12731] = !f[237] && !f[261] && f[239] && !f[215];
	assign leaf[12732] = !f[237] && !f[261] && f[239] && f[215];
	assign leaf[12733] = !f[237] && f[261] && !f[181] && !f[265];
	assign leaf[12734] = !f[237] && f[261] && !f[181] && f[265];
	assign leaf[12735] = !f[237] && f[261] && f[181] && !f[629];
	assign leaf[12736] = !f[237] && f[261] && f[181] && f[629];
	assign leaf[12737] = f[237] && !f[261] && !f[185] && !f[271];
	assign leaf[12738] = f[237] && !f[261] && !f[185] && f[271];
	assign leaf[12739] = f[237] && !f[261] && f[185] && !f[215];
	assign leaf[12740] = f[237] && !f[261] && f[185] && f[215];
	assign leaf[12741] = f[237] && f[261] && !f[272] && !f[663];
	assign leaf[12742] = f[237] && f[261] && !f[272] && f[663];
	assign leaf[12743] = f[237] && f[261] && f[272] && !f[241];
	assign leaf[12744] = f[237] && f[261] && f[272] && f[241];
	
	// Tree 935, Classifier 5, Iteration: 93
	assign leaf[12745] = !f[276] && !f[434] && !f[520] && !f[322];
	assign leaf[12746] = !f[276] && !f[434] && !f[520] && f[322];
	assign leaf[12747] = !f[276] && !f[434] && f[520] && !f[264];
	assign leaf[12748] = !f[276] && !f[434] && f[520] && f[264];
	assign leaf[12749] = !f[276] && f[434] && !f[325] && !f[215];
	assign leaf[12750] = !f[276] && f[434] && !f[325] && f[215];
	assign leaf[12751] = !f[276] && f[434] && f[325] && !f[352];
	assign leaf[12752] = !f[276] && f[434] && f[325] && f[352];
	assign leaf[12753] = f[276] && !f[273];
	assign leaf[12754] = f[276] && f[273] && !f[262] && !f[351];
	assign leaf[12755] = f[276] && f[273] && !f[262] && f[351];
	assign leaf[12756] = f[276] && f[273] && f[262];
	
	// Tree 936, Classifier 6, Iteration: 93
	assign leaf[12757] = !f[516] && !f[486] && !f[511] && !f[485];
	assign leaf[12758] = !f[516] && !f[486] && !f[511] && f[485];
	assign leaf[12759] = !f[516] && !f[486] && f[511] && !f[349];
	assign leaf[12760] = !f[516] && !f[486] && f[511] && f[349];
	assign leaf[12761] = !f[516] && f[486] && !f[542] && !f[133];
	assign leaf[12762] = !f[516] && f[486] && !f[542] && f[133];
	assign leaf[12763] = !f[516] && f[486] && f[542] && !f[295];
	assign leaf[12764] = !f[516] && f[486] && f[542] && f[295];
	assign leaf[12765] = f[516] && !f[432] && !f[515] && !f[380];
	assign leaf[12766] = f[516] && !f[432] && !f[515] && f[380];
	assign leaf[12767] = f[516] && !f[432] && f[515] && !f[462];
	assign leaf[12768] = f[516] && !f[432] && f[515] && f[462];
	assign leaf[12769] = f[516] && f[432] && !f[155] && !f[209];
	assign leaf[12770] = f[516] && f[432] && !f[155] && f[209];
	assign leaf[12771] = f[516] && f[432] && f[155] && !f[573];
	assign leaf[12772] = f[516] && f[432] && f[155] && f[573];
	
	// Tree 937, Classifier 7, Iteration: 93
	assign leaf[12773] = !f[349] && !f[432] && !f[488] && !f[290];
	assign leaf[12774] = !f[349] && !f[432] && !f[488] && f[290];
	assign leaf[12775] = !f[349] && !f[432] && f[488] && !f[429];
	assign leaf[12776] = !f[349] && !f[432] && f[488] && f[429];
	assign leaf[12777] = !f[349] && f[432] && !f[319] && !f[463];
	assign leaf[12778] = !f[349] && f[432] && !f[319] && f[463];
	assign leaf[12779] = !f[349] && f[432] && f[319] && !f[286];
	assign leaf[12780] = !f[349] && f[432] && f[319] && f[286];
	assign leaf[12781] = f[349] && !f[234] && !f[264] && !f[570];
	assign leaf[12782] = f[349] && !f[234] && !f[264] && f[570];
	assign leaf[12783] = f[349] && !f[234] && f[264] && !f[430];
	assign leaf[12784] = f[349] && !f[234] && f[264] && f[430];
	assign leaf[12785] = f[349] && f[234] && !f[265] && !f[405];
	assign leaf[12786] = f[349] && f[234] && !f[265] && f[405];
	assign leaf[12787] = f[349] && f[234] && f[265] && !f[289];
	assign leaf[12788] = f[349] && f[234] && f[265] && f[289];
	
	// Tree 938, Classifier 8, Iteration: 93
	assign leaf[12789] = !f[341] && !f[214] && !f[601] && !f[656];
	assign leaf[12790] = !f[341] && !f[214] && !f[601] && f[656];
	assign leaf[12791] = !f[341] && !f[214] && f[601] && !f[656];
	assign leaf[12792] = !f[341] && !f[214] && f[601] && f[656];
	assign leaf[12793] = !f[341] && f[214] && !f[573] && !f[546];
	assign leaf[12794] = !f[341] && f[214] && !f[573] && f[546];
	assign leaf[12795] = !f[341] && f[214] && f[573] && !f[435];
	assign leaf[12796] = !f[341] && f[214] && f[573] && f[435];
	assign leaf[12797] = f[341] && !f[522] && !f[466] && !f[211];
	assign leaf[12798] = f[341] && !f[522] && !f[466] && f[211];
	assign leaf[12799] = f[341] && !f[522] && f[466];
	assign leaf[12800] = f[341] && f[522] && !f[628];
	assign leaf[12801] = f[341] && f[522] && f[628];
	
	// Tree 939, Classifier 9, Iteration: 93
	assign leaf[12802] = !f[201] && !f[575] && !f[685] && !f[349];
	assign leaf[12803] = !f[201] && !f[575] && !f[685] && f[349];
	assign leaf[12804] = !f[201] && !f[575] && f[685] && !f[294];
	assign leaf[12805] = !f[201] && !f[575] && f[685] && f[294];
	assign leaf[12806] = !f[201] && f[575] && !f[518] && !f[459];
	assign leaf[12807] = !f[201] && f[575] && !f[518] && f[459];
	assign leaf[12808] = !f[201] && f[575] && f[518] && !f[179];
	assign leaf[12809] = !f[201] && f[575] && f[518] && f[179];
	assign leaf[12810] = f[201];
	
	// Tree 940, Classifier 0, Iteration: 94
	assign leaf[12811] = !f[434] && !f[526] && !f[319] && !f[291];
	assign leaf[12812] = !f[434] && !f[526] && !f[319] && f[291];
	assign leaf[12813] = !f[434] && !f[526] && f[319] && !f[468];
	assign leaf[12814] = !f[434] && !f[526] && f[319] && f[468];
	assign leaf[12815] = !f[434] && f[526] && !f[427] && !f[413];
	assign leaf[12816] = !f[434] && f[526] && !f[427] && f[413];
	assign leaf[12817] = !f[434] && f[526] && f[427] && !f[208];
	assign leaf[12818] = !f[434] && f[526] && f[427] && f[208];
	assign leaf[12819] = f[434] && !f[273] && !f[316];
	assign leaf[12820] = f[434] && !f[273] && f[316];
	assign leaf[12821] = f[434] && f[273] && !f[349];
	assign leaf[12822] = f[434] && f[273] && f[349] && !f[595];
	assign leaf[12823] = f[434] && f[273] && f[349] && f[595];
	
	// Tree 941, Classifier 1, Iteration: 94
	assign leaf[12824] = !f[490] && !f[378] && !f[322] && !f[434];
	assign leaf[12825] = !f[490] && !f[378] && !f[322] && f[434];
	assign leaf[12826] = !f[490] && !f[378] && f[322];
	assign leaf[12827] = !f[490] && f[378] && !f[630] && !f[569];
	assign leaf[12828] = !f[490] && f[378] && !f[630] && f[569];
	assign leaf[12829] = !f[490] && f[378] && f[630] && !f[407];
	assign leaf[12830] = !f[490] && f[378] && f[630] && f[407];
	assign leaf[12831] = f[490] && !f[603] && !f[516] && !f[635];
	assign leaf[12832] = f[490] && !f[603] && !f[516] && f[635];
	assign leaf[12833] = f[490] && !f[603] && f[516] && !f[236];
	assign leaf[12834] = f[490] && !f[603] && f[516] && f[236];
	assign leaf[12835] = f[490] && f[603] && !f[573] && !f[488];
	assign leaf[12836] = f[490] && f[603] && !f[573] && f[488];
	assign leaf[12837] = f[490] && f[603] && f[573] && !f[177];
	assign leaf[12838] = f[490] && f[603] && f[573] && f[177];
	
	// Tree 942, Classifier 2, Iteration: 94
	assign leaf[12839] = !f[397] && !f[154] && !f[374] && !f[493];
	assign leaf[12840] = !f[397] && !f[154] && !f[374] && f[493];
	assign leaf[12841] = !f[397] && !f[154] && f[374] && !f[182];
	assign leaf[12842] = !f[397] && !f[154] && f[374] && f[182];
	assign leaf[12843] = !f[397] && f[154] && !f[628] && !f[432];
	assign leaf[12844] = !f[397] && f[154] && !f[628] && f[432];
	assign leaf[12845] = !f[397] && f[154] && f[628] && !f[266];
	assign leaf[12846] = !f[397] && f[154] && f[628] && f[266];
	assign leaf[12847] = f[397] && !f[426] && !f[435];
	assign leaf[12848] = f[397] && !f[426] && f[435];
	assign leaf[12849] = f[397] && f[426] && !f[375];
	assign leaf[12850] = f[397] && f[426] && f[375];
	
	// Tree 943, Classifier 3, Iteration: 94
	assign leaf[12851] = !f[406] && !f[517] && !f[325] && !f[217];
	assign leaf[12852] = !f[406] && !f[517] && !f[325] && f[217];
	assign leaf[12853] = !f[406] && !f[517] && f[325] && !f[437];
	assign leaf[12854] = !f[406] && !f[517] && f[325] && f[437];
	assign leaf[12855] = !f[406] && f[517] && !f[212] && !f[178];
	assign leaf[12856] = !f[406] && f[517] && !f[212] && f[178];
	assign leaf[12857] = !f[406] && f[517] && f[212] && !f[233];
	assign leaf[12858] = !f[406] && f[517] && f[212] && f[233];
	assign leaf[12859] = f[406] && !f[466] && !f[300] && !f[544];
	assign leaf[12860] = f[406] && !f[466] && !f[300] && f[544];
	assign leaf[12861] = f[406] && !f[466] && f[300] && !f[574];
	assign leaf[12862] = f[406] && !f[466] && f[300] && f[574];
	assign leaf[12863] = f[406] && f[466] && !f[347] && !f[291];
	assign leaf[12864] = f[406] && f[466] && !f[347] && f[291];
	assign leaf[12865] = f[406] && f[466] && f[347] && !f[318];
	assign leaf[12866] = f[406] && f[466] && f[347] && f[318];
	
	// Tree 944, Classifier 4, Iteration: 94
	assign leaf[12867] = !f[234] && !f[178] && !f[232] && !f[180];
	assign leaf[12868] = !f[234] && !f[178] && !f[232] && f[180];
	assign leaf[12869] = !f[234] && !f[178] && f[232] && !f[544];
	assign leaf[12870] = !f[234] && !f[178] && f[232] && f[544];
	assign leaf[12871] = !f[234] && f[178] && !f[179];
	assign leaf[12872] = !f[234] && f[178] && f[179] && !f[352];
	assign leaf[12873] = !f[234] && f[178] && f[179] && f[352];
	assign leaf[12874] = f[234] && !f[290] && !f[273] && !f[150];
	assign leaf[12875] = f[234] && !f[290] && !f[273] && f[150];
	assign leaf[12876] = f[234] && !f[290] && f[273];
	assign leaf[12877] = f[234] && f[290] && !f[209] && !f[239];
	assign leaf[12878] = f[234] && f[290] && !f[209] && f[239];
	assign leaf[12879] = f[234] && f[290] && f[209] && !f[239];
	assign leaf[12880] = f[234] && f[290] && f[209] && f[239];
	
	// Tree 945, Classifier 5, Iteration: 94
	assign leaf[12881] = !f[612] && !f[147] && !f[258] && !f[155];
	assign leaf[12882] = !f[612] && !f[147] && !f[258] && f[155];
	assign leaf[12883] = !f[612] && !f[147] && f[258] && !f[399];
	assign leaf[12884] = !f[612] && !f[147] && f[258] && f[399];
	assign leaf[12885] = !f[612] && f[147] && !f[204] && !f[208];
	assign leaf[12886] = !f[612] && f[147] && !f[204] && f[208];
	assign leaf[12887] = !f[612] && f[147] && f[204] && !f[498];
	assign leaf[12888] = !f[612] && f[147] && f[204] && f[498];
	assign leaf[12889] = f[612];
	
	// Tree 946, Classifier 6, Iteration: 94
	assign leaf[12890] = !f[656] && !f[146] && !f[351] && !f[299];
	assign leaf[12891] = !f[656] && !f[146] && !f[351] && f[299];
	assign leaf[12892] = !f[656] && !f[146] && f[351] && !f[491];
	assign leaf[12893] = !f[656] && !f[146] && f[351] && f[491];
	assign leaf[12894] = !f[656] && f[146];
	assign leaf[12895] = f[656] && !f[181] && !f[157] && !f[266];
	assign leaf[12896] = f[656] && !f[181] && !f[157] && f[266];
	assign leaf[12897] = f[656] && !f[181] && f[157] && !f[242];
	assign leaf[12898] = f[656] && !f[181] && f[157] && f[242];
	assign leaf[12899] = f[656] && f[181] && !f[605];
	assign leaf[12900] = f[656] && f[181] && f[605] && !f[578];
	assign leaf[12901] = f[656] && f[181] && f[605] && f[578];
	
	// Tree 947, Classifier 7, Iteration: 94
	assign leaf[12902] = !f[605] && !f[472] && !f[482] && !f[411];
	assign leaf[12903] = !f[605] && !f[472] && !f[482] && f[411];
	assign leaf[12904] = !f[605] && !f[472] && f[482] && !f[429];
	assign leaf[12905] = !f[605] && !f[472] && f[482] && f[429];
	assign leaf[12906] = !f[605] && f[472] && !f[431];
	assign leaf[12907] = !f[605] && f[472] && f[431];
	assign leaf[12908] = f[605] && !f[516] && !f[682] && !f[627];
	assign leaf[12909] = f[605] && !f[516] && !f[682] && f[627];
	assign leaf[12910] = f[605] && !f[516] && f[682];
	assign leaf[12911] = f[605] && f[516] && !f[524] && !f[216];
	assign leaf[12912] = f[605] && f[516] && !f[524] && f[216];
	assign leaf[12913] = f[605] && f[516] && f[524] && !f[688];
	assign leaf[12914] = f[605] && f[516] && f[524] && f[688];
	
	// Tree 948, Classifier 8, Iteration: 94
	assign leaf[12915] = !f[657] && !f[629] && !f[381] && !f[317];
	assign leaf[12916] = !f[657] && !f[629] && !f[381] && f[317];
	assign leaf[12917] = !f[657] && !f[629] && f[381] && !f[433];
	assign leaf[12918] = !f[657] && !f[629] && f[381] && f[433];
	assign leaf[12919] = !f[657] && f[629] && !f[656] && !f[461];
	assign leaf[12920] = !f[657] && f[629] && !f[656] && f[461];
	assign leaf[12921] = !f[657] && f[629] && f[656] && !f[492];
	assign leaf[12922] = !f[657] && f[629] && f[656] && f[492];
	assign leaf[12923] = f[657] && !f[630] && !f[433] && !f[346];
	assign leaf[12924] = f[657] && !f[630] && !f[433] && f[346];
	assign leaf[12925] = f[657] && !f[630] && f[433] && !f[155];
	assign leaf[12926] = f[657] && !f[630] && f[433] && f[155];
	assign leaf[12927] = f[657] && f[630] && !f[633] && !f[543];
	assign leaf[12928] = f[657] && f[630] && !f[633] && f[543];
	assign leaf[12929] = f[657] && f[630] && f[633] && !f[349];
	assign leaf[12930] = f[657] && f[630] && f[633] && f[349];
	
	// Tree 949, Classifier 9, Iteration: 94
	assign leaf[12931] = !f[536] && !f[201] && !f[599] && !f[654];
	assign leaf[12932] = !f[536] && !f[201] && !f[599] && f[654];
	assign leaf[12933] = !f[536] && !f[201] && f[599] && !f[487];
	assign leaf[12934] = !f[536] && !f[201] && f[599] && f[487];
	assign leaf[12935] = !f[536] && f[201];
	assign leaf[12936] = f[536];
	
	// Tree 950, Classifier 0, Iteration: 95
	assign leaf[12937] = !f[408] && !f[574] && !f[233] && !f[541];
	assign leaf[12938] = !f[408] && !f[574] && !f[233] && f[541];
	assign leaf[12939] = !f[408] && !f[574] && f[233] && !f[347];
	assign leaf[12940] = !f[408] && !f[574] && f[233] && f[347];
	assign leaf[12941] = !f[408] && f[574] && !f[354] && !f[190];
	assign leaf[12942] = !f[408] && f[574] && !f[354] && f[190];
	assign leaf[12943] = !f[408] && f[574] && f[354] && !f[240];
	assign leaf[12944] = !f[408] && f[574] && f[354] && f[240];
	assign leaf[12945] = f[408] && !f[464] && !f[600];
	assign leaf[12946] = f[408] && !f[464] && f[600];
	assign leaf[12947] = f[408] && f[464] && !f[571];
	assign leaf[12948] = f[408] && f[464] && f[571] && !f[577];
	assign leaf[12949] = f[408] && f[464] && f[571] && f[577];
	
	// Tree 951, Classifier 1, Iteration: 95
	assign leaf[12950] = !f[378] && !f[682] && !f[624] && !f[321];
	assign leaf[12951] = !f[378] && !f[682] && !f[624] && f[321];
	assign leaf[12952] = !f[378] && !f[682] && f[624] && !f[379];
	assign leaf[12953] = !f[378] && !f[682] && f[624] && f[379];
	assign leaf[12954] = !f[378] && f[682];
	assign leaf[12955] = f[378] && !f[294] && !f[539] && !f[403];
	assign leaf[12956] = f[378] && !f[294] && !f[539] && f[403];
	assign leaf[12957] = f[378] && !f[294] && f[539];
	assign leaf[12958] = f[378] && f[294] && !f[322];
	assign leaf[12959] = f[378] && f[294] && f[322] && !f[177];
	assign leaf[12960] = f[378] && f[294] && f[322] && f[177];
	
	// Tree 952, Classifier 2, Iteration: 95
	assign leaf[12961] = !f[513] && !f[259] && !f[580] && !f[662];
	assign leaf[12962] = !f[513] && !f[259] && !f[580] && f[662];
	assign leaf[12963] = !f[513] && !f[259] && f[580] && !f[497];
	assign leaf[12964] = !f[513] && !f[259] && f[580] && f[497];
	assign leaf[12965] = !f[513] && f[259] && !f[579] && !f[428];
	assign leaf[12966] = !f[513] && f[259] && !f[579] && f[428];
	assign leaf[12967] = !f[513] && f[259] && f[579] && !f[293];
	assign leaf[12968] = !f[513] && f[259] && f[579] && f[293];
	assign leaf[12969] = f[513] && !f[287] && !f[295] && !f[317];
	assign leaf[12970] = f[513] && !f[287] && !f[295] && f[317];
	assign leaf[12971] = f[513] && !f[287] && f[295] && !f[431];
	assign leaf[12972] = f[513] && !f[287] && f[295] && f[431];
	assign leaf[12973] = f[513] && f[287] && !f[595] && !f[579];
	assign leaf[12974] = f[513] && f[287] && !f[595] && f[579];
	assign leaf[12975] = f[513] && f[287] && f[595];
	
	// Tree 953, Classifier 3, Iteration: 95
	assign leaf[12976] = !f[401] && !f[347] && !f[321] && !f[570];
	assign leaf[12977] = !f[401] && !f[347] && !f[321] && f[570];
	assign leaf[12978] = !f[401] && !f[347] && f[321] && !f[127];
	assign leaf[12979] = !f[401] && !f[347] && f[321] && f[127];
	assign leaf[12980] = !f[401] && f[347] && !f[321] && !f[174];
	assign leaf[12981] = !f[401] && f[347] && !f[321] && f[174];
	assign leaf[12982] = !f[401] && f[347] && f[321] && !f[430];
	assign leaf[12983] = !f[401] && f[347] && f[321] && f[430];
	assign leaf[12984] = f[401] && !f[651] && !f[384] && !f[328];
	assign leaf[12985] = f[401] && !f[651] && !f[384] && f[328];
	assign leaf[12986] = f[401] && !f[651] && f[384] && !f[292];
	assign leaf[12987] = f[401] && !f[651] && f[384] && f[292];
	assign leaf[12988] = f[401] && f[651] && !f[565] && !f[568];
	assign leaf[12989] = f[401] && f[651] && !f[565] && f[568];
	assign leaf[12990] = f[401] && f[651] && f[565] && !f[455];
	assign leaf[12991] = f[401] && f[651] && f[565] && f[455];
	
	// Tree 954, Classifier 4, Iteration: 95
	assign leaf[12992] = !f[741] && !f[97] && !f[381] && !f[379];
	assign leaf[12993] = !f[741] && !f[97] && !f[381] && f[379];
	assign leaf[12994] = !f[741] && !f[97] && f[381] && !f[373];
	assign leaf[12995] = !f[741] && !f[97] && f[381] && f[373];
	assign leaf[12996] = !f[741] && f[97];
	assign leaf[12997] = f[741] && !f[462];
	assign leaf[12998] = f[741] && f[462];
	
	// Tree 955, Classifier 5, Iteration: 95
	assign leaf[12999] = !f[636] && !f[177] && !f[315] && !f[232];
	assign leaf[13000] = !f[636] && !f[177] && !f[315] && f[232];
	assign leaf[13001] = !f[636] && !f[177] && f[315] && !f[204];
	assign leaf[13002] = !f[636] && !f[177] && f[315] && f[204];
	assign leaf[13003] = !f[636] && f[177] && !f[128] && !f[206];
	assign leaf[13004] = !f[636] && f[177] && !f[128] && f[206];
	assign leaf[13005] = !f[636] && f[177] && f[128] && !f[261];
	assign leaf[13006] = !f[636] && f[177] && f[128] && f[261];
	assign leaf[13007] = f[636] && !f[344] && !f[406] && !f[266];
	assign leaf[13008] = f[636] && !f[344] && !f[406] && f[266];
	assign leaf[13009] = f[636] && !f[344] && f[406] && !f[598];
	assign leaf[13010] = f[636] && !f[344] && f[406] && f[598];
	assign leaf[13011] = f[636] && f[344] && !f[260] && !f[378];
	assign leaf[13012] = f[636] && f[344] && !f[260] && f[378];
	assign leaf[13013] = f[636] && f[344] && f[260] && !f[660];
	assign leaf[13014] = f[636] && f[344] && f[260] && f[660];
	
	// Tree 956, Classifier 6, Iteration: 95
	assign leaf[13015] = !f[661] && !f[262] && !f[521] && !f[490];
	assign leaf[13016] = !f[661] && !f[262] && !f[521] && f[490];
	assign leaf[13017] = !f[661] && !f[262] && f[521] && !f[348];
	assign leaf[13018] = !f[661] && !f[262] && f[521] && f[348];
	assign leaf[13019] = !f[661] && f[262] && !f[124] && !f[568];
	assign leaf[13020] = !f[661] && f[262] && !f[124] && f[568];
	assign leaf[13021] = !f[661] && f[262] && f[124] && !f[156];
	assign leaf[13022] = !f[661] && f[262] && f[124] && f[156];
	assign leaf[13023] = f[661] && !f[552] && !f[321] && !f[237];
	assign leaf[13024] = f[661] && !f[552] && !f[321] && f[237];
	assign leaf[13025] = f[661] && !f[552] && f[321];
	assign leaf[13026] = f[661] && f[552] && !f[233] && !f[234];
	assign leaf[13027] = f[661] && f[552] && !f[233] && f[234];
	assign leaf[13028] = f[661] && f[552] && f[233] && !f[128];
	assign leaf[13029] = f[661] && f[552] && f[233] && f[128];
	
	// Tree 957, Classifier 7, Iteration: 95
	assign leaf[13030] = !f[241] && !f[350] && !f[434] && !f[349];
	assign leaf[13031] = !f[241] && !f[350] && !f[434] && f[349];
	assign leaf[13032] = !f[241] && !f[350] && f[434] && !f[653];
	assign leaf[13033] = !f[241] && !f[350] && f[434] && f[653];
	assign leaf[13034] = !f[241] && f[350] && !f[329] && !f[430];
	assign leaf[13035] = !f[241] && f[350] && !f[329] && f[430];
	assign leaf[13036] = !f[241] && f[350] && f[329] && !f[657];
	assign leaf[13037] = !f[241] && f[350] && f[329] && f[657];
	assign leaf[13038] = f[241] && !f[229] && !f[356] && !f[322];
	assign leaf[13039] = f[241] && !f[229] && !f[356] && f[322];
	assign leaf[13040] = f[241] && !f[229] && f[356] && !f[245];
	assign leaf[13041] = f[241] && !f[229] && f[356] && f[245];
	assign leaf[13042] = f[241] && f[229] && !f[541] && !f[627];
	assign leaf[13043] = f[241] && f[229] && !f[541] && f[627];
	assign leaf[13044] = f[241] && f[229] && f[541];
	
	// Tree 958, Classifier 8, Iteration: 95
	assign leaf[13045] = !f[571] && !f[595] && !f[569] && !f[513];
	assign leaf[13046] = !f[571] && !f[595] && !f[569] && f[513];
	assign leaf[13047] = !f[571] && !f[595] && f[569] && !f[494];
	assign leaf[13048] = !f[571] && !f[595] && f[569] && f[494];
	assign leaf[13049] = !f[571] && f[595] && !f[456] && !f[605];
	assign leaf[13050] = !f[571] && f[595] && !f[456] && f[605];
	assign leaf[13051] = !f[571] && f[595] && f[456] && !f[325];
	assign leaf[13052] = !f[571] && f[595] && f[456] && f[325];
	assign leaf[13053] = f[571] && !f[680] && !f[569] && !f[216];
	assign leaf[13054] = f[571] && !f[680] && !f[569] && f[216];
	assign leaf[13055] = f[571] && !f[680] && f[569] && !f[158];
	assign leaf[13056] = f[571] && !f[680] && f[569] && f[158];
	assign leaf[13057] = f[571] && f[680] && !f[683] && !f[541];
	assign leaf[13058] = f[571] && f[680] && !f[683] && f[541];
	assign leaf[13059] = f[571] && f[680] && f[683] && !f[569];
	assign leaf[13060] = f[571] && f[680] && f[683] && f[569];
	
	// Tree 959, Classifier 9, Iteration: 95
	assign leaf[13061] = !f[174] && !f[322] && !f[402] && !f[456];
	assign leaf[13062] = !f[174] && !f[322] && !f[402] && f[456];
	assign leaf[13063] = !f[174] && !f[322] && f[402] && !f[455];
	assign leaf[13064] = !f[174] && !f[322] && f[402] && f[455];
	assign leaf[13065] = !f[174] && f[322] && !f[157] && !f[540];
	assign leaf[13066] = !f[174] && f[322] && !f[157] && f[540];
	assign leaf[13067] = !f[174] && f[322] && f[157] && !f[315];
	assign leaf[13068] = !f[174] && f[322] && f[157] && f[315];
	assign leaf[13069] = f[174];
	
	// Tree 960, Classifier 0, Iteration: 96
	assign leaf[13070] = !f[294] && !f[547] && !f[659] && !f[550];
	assign leaf[13071] = !f[294] && !f[547] && !f[659] && f[550];
	assign leaf[13072] = !f[294] && !f[547] && f[659] && !f[432];
	assign leaf[13073] = !f[294] && !f[547] && f[659] && f[432];
	assign leaf[13074] = !f[294] && f[547] && !f[660] && !f[599];
	assign leaf[13075] = !f[294] && f[547] && !f[660] && f[599];
	assign leaf[13076] = !f[294] && f[547] && f[660];
	assign leaf[13077] = f[294] && !f[435] && !f[331] && !f[327];
	assign leaf[13078] = f[294] && !f[435] && !f[331] && f[327];
	assign leaf[13079] = f[294] && !f[435] && f[331] && !f[539];
	assign leaf[13080] = f[294] && !f[435] && f[331] && f[539];
	assign leaf[13081] = f[294] && f[435] && !f[434] && !f[244];
	assign leaf[13082] = f[294] && f[435] && !f[434] && f[244];
	assign leaf[13083] = f[294] && f[435] && f[434] && !f[130];
	assign leaf[13084] = f[294] && f[435] && f[434] && f[130];
	
	// Tree 961, Classifier 1, Iteration: 96
	assign leaf[13085] = !f[265] && !f[155] && !f[241] && !f[295];
	assign leaf[13086] = !f[265] && !f[155] && !f[241] && f[295];
	assign leaf[13087] = !f[265] && !f[155] && f[241] && !f[324];
	assign leaf[13088] = !f[265] && !f[155] && f[241] && f[324];
	assign leaf[13089] = !f[265] && f[155] && !f[239] && !f[406];
	assign leaf[13090] = !f[265] && f[155] && !f[239] && f[406];
	assign leaf[13091] = !f[265] && f[155] && f[239] && !f[487];
	assign leaf[13092] = !f[265] && f[155] && f[239] && f[487];
	assign leaf[13093] = f[265] && !f[159] && !f[349] && !f[157];
	assign leaf[13094] = f[265] && !f[159] && !f[349] && f[157];
	assign leaf[13095] = f[265] && !f[159] && f[349] && !f[431];
	assign leaf[13096] = f[265] && !f[159] && f[349] && f[431];
	assign leaf[13097] = f[265] && f[159] && !f[406];
	assign leaf[13098] = f[265] && f[159] && f[406] && !f[486];
	assign leaf[13099] = f[265] && f[159] && f[406] && f[486];
	
	// Tree 962, Classifier 2, Iteration: 96
	assign leaf[13100] = !f[715] && !f[121] && !f[570] && !f[296];
	assign leaf[13101] = !f[715] && !f[121] && !f[570] && f[296];
	assign leaf[13102] = !f[715] && !f[121] && f[570] && !f[400];
	assign leaf[13103] = !f[715] && !f[121] && f[570] && f[400];
	assign leaf[13104] = !f[715] && f[121] && !f[232] && !f[128];
	assign leaf[13105] = !f[715] && f[121] && !f[232] && f[128];
	assign leaf[13106] = !f[715] && f[121] && f[232];
	assign leaf[13107] = f[715] && !f[494] && !f[178];
	assign leaf[13108] = f[715] && !f[494] && f[178];
	assign leaf[13109] = f[715] && f[494];
	
	// Tree 963, Classifier 3, Iteration: 96
	assign leaf[13110] = !f[427] && !f[241] && !f[719] && !f[518];
	assign leaf[13111] = !f[427] && !f[241] && !f[719] && f[518];
	assign leaf[13112] = !f[427] && !f[241] && f[719];
	assign leaf[13113] = !f[427] && f[241] && !f[303] && !f[184];
	assign leaf[13114] = !f[427] && f[241] && !f[303] && f[184];
	assign leaf[13115] = !f[427] && f[241] && f[303] && !f[235];
	assign leaf[13116] = !f[427] && f[241] && f[303] && f[235];
	assign leaf[13117] = f[427] && !f[437] && !f[236] && !f[327];
	assign leaf[13118] = f[427] && !f[437] && !f[236] && f[327];
	assign leaf[13119] = f[427] && !f[437] && f[236] && !f[215];
	assign leaf[13120] = f[427] && !f[437] && f[236] && f[215];
	assign leaf[13121] = f[427] && f[437] && !f[428];
	assign leaf[13122] = f[427] && f[437] && f[428] && !f[241];
	assign leaf[13123] = f[427] && f[437] && f[428] && f[241];
	
	// Tree 964, Classifier 4, Iteration: 96
	assign leaf[13124] = !f[400] && !f[349] && !f[211] && !f[294];
	assign leaf[13125] = !f[400] && !f[349] && !f[211] && f[294];
	assign leaf[13126] = !f[400] && !f[349] && f[211] && !f[237];
	assign leaf[13127] = !f[400] && !f[349] && f[211] && f[237];
	assign leaf[13128] = !f[400] && f[349] && !f[179] && !f[319];
	assign leaf[13129] = !f[400] && f[349] && !f[179] && f[319];
	assign leaf[13130] = !f[400] && f[349] && f[179] && !f[206];
	assign leaf[13131] = !f[400] && f[349] && f[179] && f[206];
	assign leaf[13132] = f[400] && !f[457] && !f[628] && !f[213];
	assign leaf[13133] = f[400] && !f[457] && !f[628] && f[213];
	assign leaf[13134] = f[400] && !f[457] && f[628] && !f[517];
	assign leaf[13135] = f[400] && !f[457] && f[628] && f[517];
	assign leaf[13136] = f[400] && f[457] && !f[439] && !f[437];
	assign leaf[13137] = f[400] && f[457] && !f[439] && f[437];
	assign leaf[13138] = f[400] && f[457] && f[439] && !f[520];
	assign leaf[13139] = f[400] && f[457] && f[439] && f[520];
	
	// Tree 965, Classifier 5, Iteration: 96
	assign leaf[13140] = !f[380] && !f[686] && !f[549] && !f[293];
	assign leaf[13141] = !f[380] && !f[686] && !f[549] && f[293];
	assign leaf[13142] = !f[380] && !f[686] && f[549] && !f[427];
	assign leaf[13143] = !f[380] && !f[686] && f[549] && f[427];
	assign leaf[13144] = !f[380] && f[686] && !f[289] && !f[296];
	assign leaf[13145] = !f[380] && f[686] && !f[289] && f[296];
	assign leaf[13146] = !f[380] && f[686] && f[289] && !f[572];
	assign leaf[13147] = !f[380] && f[686] && f[289] && f[572];
	assign leaf[13148] = f[380] && !f[248] && !f[342] && !f[522];
	assign leaf[13149] = f[380] && !f[248] && !f[342] && f[522];
	assign leaf[13150] = f[380] && !f[248] && f[342] && !f[347];
	assign leaf[13151] = f[380] && !f[248] && f[342] && f[347];
	assign leaf[13152] = f[380] && f[248] && !f[219];
	assign leaf[13153] = f[380] && f[248] && f[219];
	
	// Tree 966, Classifier 6, Iteration: 96
	assign leaf[13154] = !f[267] && !f[120] && !f[237] && !f[155];
	assign leaf[13155] = !f[267] && !f[120] && !f[237] && f[155];
	assign leaf[13156] = !f[267] && !f[120] && f[237] && !f[634];
	assign leaf[13157] = !f[267] && !f[120] && f[237] && f[634];
	assign leaf[13158] = !f[267] && f[120];
	assign leaf[13159] = f[267] && !f[321] && !f[659] && !f[551];
	assign leaf[13160] = f[267] && !f[321] && !f[659] && f[551];
	assign leaf[13161] = f[267] && !f[321] && f[659];
	assign leaf[13162] = f[267] && f[321] && !f[181] && !f[433];
	assign leaf[13163] = f[267] && f[321] && !f[181] && f[433];
	assign leaf[13164] = f[267] && f[321] && f[181] && !f[495];
	assign leaf[13165] = f[267] && f[321] && f[181] && f[495];
	
	// Tree 967, Classifier 7, Iteration: 96
	assign leaf[13166] = !f[472] && !f[202] && !f[262] && !f[292];
	assign leaf[13167] = !f[472] && !f[202] && !f[262] && f[292];
	assign leaf[13168] = !f[472] && !f[202] && f[262] && !f[265];
	assign leaf[13169] = !f[472] && !f[202] && f[262] && f[265];
	assign leaf[13170] = !f[472] && f[202] && !f[568] && !f[598];
	assign leaf[13171] = !f[472] && f[202] && !f[568] && f[598];
	assign leaf[13172] = !f[472] && f[202] && f[568];
	assign leaf[13173] = f[472] && !f[457];
	assign leaf[13174] = f[472] && f[457];
	
	// Tree 968, Classifier 8, Iteration: 96
	assign leaf[13175] = !f[442] && !f[258] && !f[526] && !f[601];
	assign leaf[13176] = !f[442] && !f[258] && !f[526] && f[601];
	assign leaf[13177] = !f[442] && !f[258] && f[526] && !f[484];
	assign leaf[13178] = !f[442] && !f[258] && f[526] && f[484];
	assign leaf[13179] = !f[442] && f[258] && !f[682] && !f[633];
	assign leaf[13180] = !f[442] && f[258] && !f[682] && f[633];
	assign leaf[13181] = !f[442] && f[258] && f[682];
	assign leaf[13182] = f[442] && !f[291] && !f[211];
	assign leaf[13183] = f[442] && !f[291] && f[211] && !f[598];
	assign leaf[13184] = f[442] && !f[291] && f[211] && f[598];
	assign leaf[13185] = f[442] && f[291] && !f[386];
	assign leaf[13186] = f[442] && f[291] && f[386];
	
	// Tree 969, Classifier 9, Iteration: 96
	assign leaf[13187] = !f[408] && !f[468] && !f[157] && !f[410];
	assign leaf[13188] = !f[408] && !f[468] && !f[157] && f[410];
	assign leaf[13189] = !f[408] && !f[468] && f[157] && !f[521];
	assign leaf[13190] = !f[408] && !f[468] && f[157] && f[521];
	assign leaf[13191] = !f[408] && f[468] && !f[517] && !f[574];
	assign leaf[13192] = !f[408] && f[468] && !f[517] && f[574];
	assign leaf[13193] = !f[408] && f[468] && f[517] && !f[470];
	assign leaf[13194] = !f[408] && f[468] && f[517] && f[470];
	assign leaf[13195] = f[408] && !f[467] && !f[412] && !f[352];
	assign leaf[13196] = f[408] && !f[467] && !f[412] && f[352];
	assign leaf[13197] = f[408] && !f[467] && f[412] && !f[328];
	assign leaf[13198] = f[408] && !f[467] && f[412] && f[328];
	assign leaf[13199] = f[408] && f[467] && !f[384] && !f[635];
	assign leaf[13200] = f[408] && f[467] && !f[384] && f[635];
	assign leaf[13201] = f[408] && f[467] && f[384] && !f[322];
	assign leaf[13202] = f[408] && f[467] && f[384] && f[322];
	
	// Tree 970, Classifier 0, Iteration: 97
	assign leaf[13203] = !f[555] && !f[468] && !f[602] && !f[460];
	assign leaf[13204] = !f[555] && !f[468] && !f[602] && f[460];
	assign leaf[13205] = !f[555] && !f[468] && f[602] && !f[432];
	assign leaf[13206] = !f[555] && !f[468] && f[602] && f[432];
	assign leaf[13207] = !f[555] && f[468] && !f[295] && !f[268];
	assign leaf[13208] = !f[555] && f[468] && !f[295] && f[268];
	assign leaf[13209] = !f[555] && f[468] && f[295] && !f[569];
	assign leaf[13210] = !f[555] && f[468] && f[295] && f[569];
	assign leaf[13211] = f[555] && !f[398];
	assign leaf[13212] = f[555] && f[398];
	
	// Tree 971, Classifier 1, Iteration: 97
	assign leaf[13213] = !f[658] && !f[517] && !f[184] && !f[238];
	assign leaf[13214] = !f[658] && !f[517] && !f[184] && f[238];
	assign leaf[13215] = !f[658] && !f[517] && f[184] && !f[578];
	assign leaf[13216] = !f[658] && !f[517] && f[184] && f[578];
	assign leaf[13217] = !f[658] && f[517] && !f[241] && !f[380];
	assign leaf[13218] = !f[658] && f[517] && !f[241] && f[380];
	assign leaf[13219] = !f[658] && f[517] && f[241] && !f[349];
	assign leaf[13220] = !f[658] && f[517] && f[241] && f[349];
	assign leaf[13221] = f[658] && !f[266] && !f[181];
	assign leaf[13222] = f[658] && !f[266] && f[181] && !f[464];
	assign leaf[13223] = f[658] && !f[266] && f[181] && f[464];
	assign leaf[13224] = f[658] && f[266] && !f[517] && !f[377];
	assign leaf[13225] = f[658] && f[266] && !f[517] && f[377];
	assign leaf[13226] = f[658] && f[266] && f[517] && !f[600];
	assign leaf[13227] = f[658] && f[266] && f[517] && f[600];
	
	// Tree 972, Classifier 2, Iteration: 97
	assign leaf[13228] = !f[94] && !f[133] && !f[543] && !f[554];
	assign leaf[13229] = !f[94] && !f[133] && !f[543] && f[554];
	assign leaf[13230] = !f[94] && !f[133] && f[543] && !f[570];
	assign leaf[13231] = !f[94] && !f[133] && f[543] && f[570];
	assign leaf[13232] = !f[94] && f[133] && !f[273] && !f[574];
	assign leaf[13233] = !f[94] && f[133] && !f[273] && f[574];
	assign leaf[13234] = !f[94] && f[133] && f[273] && !f[577];
	assign leaf[13235] = !f[94] && f[133] && f[273] && f[577];
	assign leaf[13236] = f[94] && !f[149];
	assign leaf[13237] = f[94] && f[149];
	
	// Tree 973, Classifier 3, Iteration: 97
	assign leaf[13238] = !f[492] && !f[598] && !f[575] && !f[600];
	assign leaf[13239] = !f[492] && !f[598] && !f[575] && f[600];
	assign leaf[13240] = !f[492] && !f[598] && f[575] && !f[354];
	assign leaf[13241] = !f[492] && !f[598] && f[575] && f[354];
	assign leaf[13242] = !f[492] && f[598] && !f[629] && !f[495];
	assign leaf[13243] = !f[492] && f[598] && !f[629] && f[495];
	assign leaf[13244] = !f[492] && f[598] && f[629] && !f[573];
	assign leaf[13245] = !f[492] && f[598] && f[629] && f[573];
	assign leaf[13246] = f[492] && !f[468] && !f[493] && !f[293];
	assign leaf[13247] = f[492] && !f[468] && !f[493] && f[293];
	assign leaf[13248] = f[492] && !f[468] && f[493] && !f[346];
	assign leaf[13249] = f[492] && !f[468] && f[493] && f[346];
	assign leaf[13250] = f[492] && f[468] && !f[554] && !f[274];
	assign leaf[13251] = f[492] && f[468] && !f[554] && f[274];
	assign leaf[13252] = f[492] && f[468] && f[554] && !f[297];
	assign leaf[13253] = f[492] && f[468] && f[554] && f[297];
	
	// Tree 974, Classifier 4, Iteration: 97
	assign leaf[13254] = !f[708] && !f[267] && !f[184] && !f[215];
	assign leaf[13255] = !f[708] && !f[267] && !f[184] && f[215];
	assign leaf[13256] = !f[708] && !f[267] && f[184] && !f[268];
	assign leaf[13257] = !f[708] && !f[267] && f[184] && f[268];
	assign leaf[13258] = !f[708] && f[267] && !f[242] && !f[236];
	assign leaf[13259] = !f[708] && f[267] && !f[242] && f[236];
	assign leaf[13260] = !f[708] && f[267] && f[242] && !f[497];
	assign leaf[13261] = !f[708] && f[267] && f[242] && f[497];
	assign leaf[13262] = f[708] && !f[241];
	assign leaf[13263] = f[708] && f[241];
	
	// Tree 975, Classifier 5, Iteration: 97
	assign leaf[13264] = !f[707] && !f[424] && !f[508] && !f[322];
	assign leaf[13265] = !f[707] && !f[424] && !f[508] && f[322];
	assign leaf[13266] = !f[707] && !f[424] && f[508] && !f[301];
	assign leaf[13267] = !f[707] && !f[424] && f[508] && f[301];
	assign leaf[13268] = !f[707] && f[424] && !f[357];
	assign leaf[13269] = !f[707] && f[424] && f[357];
	assign leaf[13270] = f[707];
	
	// Tree 976, Classifier 6, Iteration: 97
	assign leaf[13271] = !f[547] && !f[631] && !f[603] && !f[463];
	assign leaf[13272] = !f[547] && !f[631] && !f[603] && f[463];
	assign leaf[13273] = !f[547] && !f[631] && f[603] && !f[493];
	assign leaf[13274] = !f[547] && !f[631] && f[603] && f[493];
	assign leaf[13275] = !f[547] && f[631] && !f[178] && !f[267];
	assign leaf[13276] = !f[547] && f[631] && !f[178] && f[267];
	assign leaf[13277] = !f[547] && f[631] && f[178] && !f[456];
	assign leaf[13278] = !f[547] && f[631] && f[178] && f[456];
	assign leaf[13279] = f[547] && !f[488] && !f[572] && !f[513];
	assign leaf[13280] = f[547] && !f[488] && !f[572] && f[513];
	assign leaf[13281] = f[547] && !f[488] && f[572] && !f[154];
	assign leaf[13282] = f[547] && !f[488] && f[572] && f[154];
	assign leaf[13283] = f[547] && f[488] && !f[631] && !f[514];
	assign leaf[13284] = f[547] && f[488] && !f[631] && f[514];
	assign leaf[13285] = f[547] && f[488] && f[631] && !f[573];
	assign leaf[13286] = f[547] && f[488] && f[631] && f[573];
	
	// Tree 977, Classifier 7, Iteration: 97
	assign leaf[13287] = !f[359] && !f[206] && !f[260] && !f[154];
	assign leaf[13288] = !f[359] && !f[206] && !f[260] && f[154];
	assign leaf[13289] = !f[359] && !f[206] && f[260] && !f[291];
	assign leaf[13290] = !f[359] && !f[206] && f[260] && f[291];
	assign leaf[13291] = !f[359] && f[206] && !f[327] && !f[259];
	assign leaf[13292] = !f[359] && f[206] && !f[327] && f[259];
	assign leaf[13293] = !f[359] && f[206] && f[327] && !f[520];
	assign leaf[13294] = !f[359] && f[206] && f[327] && f[520];
	assign leaf[13295] = f[359] && !f[683] && !f[427];
	assign leaf[13296] = f[359] && !f[683] && f[427];
	assign leaf[13297] = f[359] && f[683];
	
	// Tree 978, Classifier 8, Iteration: 97
	assign leaf[13298] = !f[211] && !f[636] && !f[154] && !f[569];
	assign leaf[13299] = !f[211] && !f[636] && !f[154] && f[569];
	assign leaf[13300] = !f[211] && !f[636] && f[154] && !f[322];
	assign leaf[13301] = !f[211] && !f[636] && f[154] && f[322];
	assign leaf[13302] = !f[211] && f[636] && !f[578] && !f[128];
	assign leaf[13303] = !f[211] && f[636] && !f[578] && f[128];
	assign leaf[13304] = !f[211] && f[636] && f[578] && !f[572];
	assign leaf[13305] = !f[211] && f[636] && f[578] && f[572];
	assign leaf[13306] = f[211] && !f[210] && !f[594] && !f[431];
	assign leaf[13307] = f[211] && !f[210] && !f[594] && f[431];
	assign leaf[13308] = f[211] && !f[210] && f[594] && !f[463];
	assign leaf[13309] = f[211] && !f[210] && f[594] && f[463];
	assign leaf[13310] = f[211] && f[210] && !f[263] && !f[273];
	assign leaf[13311] = f[211] && f[210] && !f[263] && f[273];
	assign leaf[13312] = f[211] && f[210] && f[263] && !f[204];
	assign leaf[13313] = f[211] && f[210] && f[263] && f[204];
	
	// Tree 979, Classifier 9, Iteration: 97
	assign leaf[13314] = !f[191] && !f[326] && !f[396] && !f[462];
	assign leaf[13315] = !f[191] && !f[326] && !f[396] && f[462];
	assign leaf[13316] = !f[191] && !f[326] && f[396] && !f[398];
	assign leaf[13317] = !f[191] && !f[326] && f[396] && f[398];
	assign leaf[13318] = !f[191] && f[326] && !f[271] && !f[330];
	assign leaf[13319] = !f[191] && f[326] && !f[271] && f[330];
	assign leaf[13320] = !f[191] && f[326] && f[271] && !f[356];
	assign leaf[13321] = !f[191] && f[326] && f[271] && f[356];
	assign leaf[13322] = f[191] && !f[188];
	assign leaf[13323] = f[191] && f[188];
	
	// Tree 980, Classifier 0, Iteration: 98
	assign leaf[13324] = !f[425] && !f[542] && !f[541] && !f[271];
	assign leaf[13325] = !f[425] && !f[542] && !f[541] && f[271];
	assign leaf[13326] = !f[425] && !f[542] && f[541] && !f[382];
	assign leaf[13327] = !f[425] && !f[542] && f[541] && f[382];
	assign leaf[13328] = !f[425] && f[542] && !f[247] && !f[510];
	assign leaf[13329] = !f[425] && f[542] && !f[247] && f[510];
	assign leaf[13330] = !f[425] && f[542] && f[247];
	assign leaf[13331] = f[425] && !f[471] && !f[396] && !f[343];
	assign leaf[13332] = f[425] && !f[471] && !f[396] && f[343];
	assign leaf[13333] = f[425] && !f[471] && f[396];
	assign leaf[13334] = f[425] && f[471] && !f[317];
	assign leaf[13335] = f[425] && f[471] && f[317];
	
	// Tree 981, Classifier 1, Iteration: 98
	assign leaf[13336] = !f[320] && !f[687] && !f[373] && !f[657];
	assign leaf[13337] = !f[320] && !f[687] && !f[373] && f[657];
	assign leaf[13338] = !f[320] && !f[687] && f[373];
	assign leaf[13339] = !f[320] && f[687] && !f[180];
	assign leaf[13340] = !f[320] && f[687] && f[180] && !f[154];
	assign leaf[13341] = !f[320] && f[687] && f[180] && f[154];
	assign leaf[13342] = f[320] && !f[662] && !f[460] && !f[547];
	assign leaf[13343] = f[320] && !f[662] && !f[460] && f[547];
	assign leaf[13344] = f[320] && !f[662] && f[460] && !f[405];
	assign leaf[13345] = f[320] && !f[662] && f[460] && f[405];
	assign leaf[13346] = f[320] && f[662] && !f[267];
	assign leaf[13347] = f[320] && f[662] && f[267];
	
	// Tree 982, Classifier 2, Iteration: 98
	assign leaf[13348] = !f[487] && !f[433] && !f[174] && !f[653];
	assign leaf[13349] = !f[487] && !f[433] && !f[174] && f[653];
	assign leaf[13350] = !f[487] && !f[433] && f[174] && !f[609];
	assign leaf[13351] = !f[487] && !f[433] && f[174] && f[609];
	assign leaf[13352] = !f[487] && f[433] && !f[484] && !f[382];
	assign leaf[13353] = !f[487] && f[433] && !f[484] && f[382];
	assign leaf[13354] = !f[487] && f[433] && f[484] && !f[294];
	assign leaf[13355] = !f[487] && f[433] && f[484] && f[294];
	assign leaf[13356] = f[487] && !f[630] && !f[547] && !f[653];
	assign leaf[13357] = f[487] && !f[630] && !f[547] && f[653];
	assign leaf[13358] = f[487] && !f[630] && f[547] && !f[690];
	assign leaf[13359] = f[487] && !f[630] && f[547] && f[690];
	assign leaf[13360] = f[487] && f[630] && !f[492] && !f[439];
	assign leaf[13361] = f[487] && f[630] && !f[492] && f[439];
	assign leaf[13362] = f[487] && f[630] && f[492] && !f[385];
	assign leaf[13363] = f[487] && f[630] && f[492] && f[385];
	
	// Tree 983, Classifier 3, Iteration: 98
	assign leaf[13364] = !f[240] && !f[189] && !f[356] && !f[129];
	assign leaf[13365] = !f[240] && !f[189] && !f[356] && f[129];
	assign leaf[13366] = !f[240] && !f[189] && f[356] && !f[155];
	assign leaf[13367] = !f[240] && !f[189] && f[356] && f[155];
	assign leaf[13368] = !f[240] && f[189] && !f[245] && !f[237];
	assign leaf[13369] = !f[240] && f[189] && !f[245] && f[237];
	assign leaf[13370] = !f[240] && f[189] && f[245] && !f[627];
	assign leaf[13371] = !f[240] && f[189] && f[245] && f[627];
	assign leaf[13372] = f[240] && !f[128] && !f[319] && !f[209];
	assign leaf[13373] = f[240] && !f[128] && !f[319] && f[209];
	assign leaf[13374] = f[240] && !f[128] && f[319] && !f[316];
	assign leaf[13375] = f[240] && !f[128] && f[319] && f[316];
	assign leaf[13376] = f[240] && f[128] && !f[293] && !f[404];
	assign leaf[13377] = f[240] && f[128] && !f[293] && f[404];
	assign leaf[13378] = f[240] && f[128] && f[293] && !f[244];
	assign leaf[13379] = f[240] && f[128] && f[293] && f[244];
	
	// Tree 984, Classifier 4, Iteration: 98
	assign leaf[13380] = !f[637] && !f[409] && !f[681] && !f[398];
	assign leaf[13381] = !f[637] && !f[409] && !f[681] && f[398];
	assign leaf[13382] = !f[637] && !f[409] && f[681];
	assign leaf[13383] = !f[637] && f[409] && !f[348] && !f[401];
	assign leaf[13384] = !f[637] && f[409] && !f[348] && f[401];
	assign leaf[13385] = !f[637] && f[409] && f[348] && !f[296];
	assign leaf[13386] = !f[637] && f[409] && f[348] && f[296];
	assign leaf[13387] = f[637] && !f[205] && !f[523];
	assign leaf[13388] = f[637] && !f[205] && f[523] && !f[435];
	assign leaf[13389] = f[637] && !f[205] && f[523] && f[435];
	assign leaf[13390] = f[637] && f[205] && !f[180];
	assign leaf[13391] = f[637] && f[205] && f[180];
	
	// Tree 985, Classifier 5, Iteration: 98
	assign leaf[13392] = !f[411] && !f[158] && !f[434] && !f[270];
	assign leaf[13393] = !f[411] && !f[158] && !f[434] && f[270];
	assign leaf[13394] = !f[411] && !f[158] && f[434] && !f[352];
	assign leaf[13395] = !f[411] && !f[158] && f[434] && f[352];
	assign leaf[13396] = !f[411] && f[158] && !f[243] && !f[245];
	assign leaf[13397] = !f[411] && f[158] && !f[243] && f[245];
	assign leaf[13398] = !f[411] && f[158] && f[243] && !f[434];
	assign leaf[13399] = !f[411] && f[158] && f[243] && f[434];
	assign leaf[13400] = f[411] && !f[300] && !f[593] && !f[131];
	assign leaf[13401] = f[411] && !f[300] && !f[593] && f[131];
	assign leaf[13402] = f[411] && !f[300] && f[593] && !f[237];
	assign leaf[13403] = f[411] && !f[300] && f[593] && f[237];
	assign leaf[13404] = f[411] && f[300] && !f[383];
	assign leaf[13405] = f[411] && f[300] && f[383] && !f[356];
	assign leaf[13406] = f[411] && f[300] && f[383] && f[356];
	
	// Tree 986, Classifier 6, Iteration: 98
	assign leaf[13407] = !f[516] && !f[405] && !f[240] && !f[123];
	assign leaf[13408] = !f[516] && !f[405] && !f[240] && f[123];
	assign leaf[13409] = !f[516] && !f[405] && f[240] && !f[433];
	assign leaf[13410] = !f[516] && !f[405] && f[240] && f[433];
	assign leaf[13411] = !f[516] && f[405] && !f[486] && !f[455];
	assign leaf[13412] = !f[516] && f[405] && !f[486] && f[455];
	assign leaf[13413] = !f[516] && f[405] && f[486] && !f[233];
	assign leaf[13414] = !f[516] && f[405] && f[486] && f[233];
	assign leaf[13415] = f[516] && !f[432] && !f[486] && !f[377];
	assign leaf[13416] = f[516] && !f[432] && !f[486] && f[377];
	assign leaf[13417] = f[516] && !f[432] && f[486] && !f[631];
	assign leaf[13418] = f[516] && !f[432] && f[486] && f[631];
	assign leaf[13419] = f[516] && f[432] && !f[434] && !f[633];
	assign leaf[13420] = f[516] && f[432] && !f[434] && f[633];
	assign leaf[13421] = f[516] && f[432] && f[434] && !f[216];
	assign leaf[13422] = f[516] && f[432] && f[434] && f[216];
	
	// Tree 987, Classifier 7, Iteration: 98
	assign leaf[13423] = !f[154] && !f[159] && !f[182] && !f[542];
	assign leaf[13424] = !f[154] && !f[159] && !f[182] && f[542];
	assign leaf[13425] = !f[154] && !f[159] && f[182] && !f[290];
	assign leaf[13426] = !f[154] && !f[159] && f[182] && f[290];
	assign leaf[13427] = !f[154] && f[159];
	assign leaf[13428] = f[154] && !f[403] && !f[186] && !f[463];
	assign leaf[13429] = f[154] && !f[403] && !f[186] && f[463];
	assign leaf[13430] = f[154] && !f[403] && f[186] && !f[233];
	assign leaf[13431] = f[154] && !f[403] && f[186] && f[233];
	assign leaf[13432] = f[154] && f[403] && !f[684];
	assign leaf[13433] = f[154] && f[403] && f[684];
	
	// Tree 988, Classifier 8, Iteration: 98
	assign leaf[13434] = !f[458] && !f[512] && !f[488] && !f[517];
	assign leaf[13435] = !f[458] && !f[512] && !f[488] && f[517];
	assign leaf[13436] = !f[458] && !f[512] && f[488] && !f[517];
	assign leaf[13437] = !f[458] && !f[512] && f[488] && f[517];
	assign leaf[13438] = !f[458] && f[512] && !f[576] && !f[348];
	assign leaf[13439] = !f[458] && f[512] && !f[576] && f[348];
	assign leaf[13440] = !f[458] && f[512] && f[576] && !f[274];
	assign leaf[13441] = !f[458] && f[512] && f[576] && f[274];
	assign leaf[13442] = f[458] && !f[489] && !f[454] && !f[294];
	assign leaf[13443] = f[458] && !f[489] && !f[454] && f[294];
	assign leaf[13444] = f[458] && !f[489] && f[454] && !f[436];
	assign leaf[13445] = f[458] && !f[489] && f[454] && f[436];
	assign leaf[13446] = f[458] && f[489] && !f[373] && !f[596];
	assign leaf[13447] = f[458] && f[489] && !f[373] && f[596];
	assign leaf[13448] = f[458] && f[489] && f[373] && !f[521];
	assign leaf[13449] = f[458] && f[489] && f[373] && f[521];
	
	// Tree 989, Classifier 9, Iteration: 98
	assign leaf[13450] = !f[186] && !f[262] && !f[205] && !f[466];
	assign leaf[13451] = !f[186] && !f[262] && !f[205] && f[466];
	assign leaf[13452] = !f[186] && !f[262] && f[205] && !f[179];
	assign leaf[13453] = !f[186] && !f[262] && f[205] && f[179];
	assign leaf[13454] = !f[186] && f[262] && !f[246] && !f[235];
	assign leaf[13455] = !f[186] && f[262] && !f[246] && f[235];
	assign leaf[13456] = !f[186] && f[262] && f[246] && !f[207];
	assign leaf[13457] = !f[186] && f[262] && f[246] && f[207];
	assign leaf[13458] = f[186] && !f[241] && !f[185] && !f[263];
	assign leaf[13459] = f[186] && !f[241] && !f[185] && f[263];
	assign leaf[13460] = f[186] && !f[241] && f[185] && !f[684];
	assign leaf[13461] = f[186] && !f[241] && f[185] && f[684];
	assign leaf[13462] = f[186] && f[241] && !f[238] && !f[183];
	assign leaf[13463] = f[186] && f[241] && !f[238] && f[183];
	assign leaf[13464] = f[186] && f[241] && f[238] && !f[491];
	assign leaf[13465] = f[186] && f[241] && f[238] && f[491];
	
	// Tree 990, Classifier 0, Iteration: 99
	assign leaf[13466] = !f[386] && !f[354] && !f[416] && !f[356];
	assign leaf[13467] = !f[386] && !f[354] && !f[416] && f[356];
	assign leaf[13468] = !f[386] && !f[354] && f[416];
	assign leaf[13469] = !f[386] && f[354] && !f[187] && !f[515];
	assign leaf[13470] = !f[386] && f[354] && !f[187] && f[515];
	assign leaf[13471] = !f[386] && f[354] && f[187] && !f[130];
	assign leaf[13472] = !f[386] && f[354] && f[187] && f[130];
	assign leaf[13473] = f[386] && !f[159] && !f[383] && !f[273];
	assign leaf[13474] = f[386] && !f[159] && !f[383] && f[273];
	assign leaf[13475] = f[386] && !f[159] && f[383] && !f[297];
	assign leaf[13476] = f[386] && !f[159] && f[383] && f[297];
	assign leaf[13477] = f[386] && f[159] && !f[570];
	assign leaf[13478] = f[386] && f[159] && f[570];
	
	// Tree 991, Classifier 1, Iteration: 99
	assign leaf[13479] = !f[708] && !f[403] && !f[714] && !f[321];
	assign leaf[13480] = !f[708] && !f[403] && !f[714] && f[321];
	assign leaf[13481] = !f[708] && !f[403] && f[714] && !f[184];
	assign leaf[13482] = !f[708] && !f[403] && f[714] && f[184];
	assign leaf[13483] = !f[708] && f[403] && !f[349];
	assign leaf[13484] = !f[708] && f[403] && f[349] && !f[155];
	assign leaf[13485] = !f[708] && f[403] && f[349] && f[155];
	assign leaf[13486] = f[708];
	
	// Tree 992, Classifier 2, Iteration: 99
	assign leaf[13487] = !f[266] && !f[317] && !f[715] && !f[513];
	assign leaf[13488] = !f[266] && !f[317] && !f[715] && f[513];
	assign leaf[13489] = !f[266] && !f[317] && f[715];
	assign leaf[13490] = !f[266] && f[317] && !f[436] && !f[566];
	assign leaf[13491] = !f[266] && f[317] && !f[436] && f[566];
	assign leaf[13492] = !f[266] && f[317] && f[436] && !f[380];
	assign leaf[13493] = !f[266] && f[317] && f[436] && f[380];
	assign leaf[13494] = f[266] && !f[542] && !f[408] && !f[488];
	assign leaf[13495] = f[266] && !f[542] && !f[408] && f[488];
	assign leaf[13496] = f[266] && !f[542] && f[408] && !f[482];
	assign leaf[13497] = f[266] && !f[542] && f[408] && f[482];
	assign leaf[13498] = f[266] && f[542] && !f[622] && !f[354];
	assign leaf[13499] = f[266] && f[542] && !f[622] && f[354];
	assign leaf[13500] = f[266] && f[542] && f[622] && !f[518];
	assign leaf[13501] = f[266] && f[542] && f[622] && f[518];
	
	// Tree 993, Classifier 3, Iteration: 99
	assign leaf[13502] = !f[411] && !f[466] && !f[179] && !f[493];
	assign leaf[13503] = !f[411] && !f[466] && !f[179] && f[493];
	assign leaf[13504] = !f[411] && !f[466] && f[179] && !f[571];
	assign leaf[13505] = !f[411] && !f[466] && f[179] && f[571];
	assign leaf[13506] = !f[411] && f[466] && !f[382] && !f[548];
	assign leaf[13507] = !f[411] && f[466] && !f[382] && f[548];
	assign leaf[13508] = !f[411] && f[466] && f[382] && !f[356];
	assign leaf[13509] = !f[411] && f[466] && f[382] && f[356];
	assign leaf[13510] = f[411] && !f[179] && !f[235] && !f[130];
	assign leaf[13511] = f[411] && !f[179] && !f[235] && f[130];
	assign leaf[13512] = f[411] && !f[179] && f[235] && !f[464];
	assign leaf[13513] = f[411] && !f[179] && f[235] && f[464];
	assign leaf[13514] = f[411] && f[179] && !f[293] && !f[264];
	assign leaf[13515] = f[411] && f[179] && !f[293] && f[264];
	assign leaf[13516] = f[411] && f[179] && f[293] && !f[234];
	assign leaf[13517] = f[411] && f[179] && f[293] && f[234];
	
	// Tree 994, Classifier 4, Iteration: 99
	assign leaf[13518] = !f[102] && !f[432] && !f[523] && !f[233];
	assign leaf[13519] = !f[102] && !f[432] && !f[523] && f[233];
	assign leaf[13520] = !f[102] && !f[432] && f[523] && !f[635];
	assign leaf[13521] = !f[102] && !f[432] && f[523] && f[635];
	assign leaf[13522] = !f[102] && f[432] && !f[511] && !f[232];
	assign leaf[13523] = !f[102] && f[432] && !f[511] && f[232];
	assign leaf[13524] = !f[102] && f[432] && f[511] && !f[515];
	assign leaf[13525] = !f[102] && f[432] && f[511] && f[515];
	assign leaf[13526] = f[102];
	
	// Tree 995, Classifier 5, Iteration: 99
	assign leaf[13527] = !f[297] && !f[215] && !f[266] && !f[127];
	assign leaf[13528] = !f[297] && !f[215] && !f[266] && f[127];
	assign leaf[13529] = !f[297] && !f[215] && f[266] && !f[623];
	assign leaf[13530] = !f[297] && !f[215] && f[266] && f[623];
	assign leaf[13531] = !f[297] && f[215] && !f[372] && !f[299];
	assign leaf[13532] = !f[297] && f[215] && !f[372] && f[299];
	assign leaf[13533] = !f[297] && f[215] && f[372] && !f[454];
	assign leaf[13534] = !f[297] && f[215] && f[372] && f[454];
	assign leaf[13535] = f[297] && !f[295] && !f[414] && !f[267];
	assign leaf[13536] = f[297] && !f[295] && !f[414] && f[267];
	assign leaf[13537] = f[297] && !f[295] && f[414];
	assign leaf[13538] = f[297] && f[295] && !f[242] && !f[342];
	assign leaf[13539] = f[297] && f[295] && !f[242] && f[342];
	assign leaf[13540] = f[297] && f[295] && f[242] && !f[156];
	assign leaf[13541] = f[297] && f[295] && f[242] && f[156];
	
	// Tree 996, Classifier 6, Iteration: 99
	assign leaf[13542] = !f[516] && !f[544] && !f[570] && !f[568];
	assign leaf[13543] = !f[516] && !f[544] && !f[570] && f[568];
	assign leaf[13544] = !f[516] && !f[544] && f[570] && !f[654];
	assign leaf[13545] = !f[516] && !f[544] && f[570] && f[654];
	assign leaf[13546] = !f[516] && f[544] && !f[457] && !f[320];
	assign leaf[13547] = !f[516] && f[544] && !f[457] && f[320];
	assign leaf[13548] = !f[516] && f[544] && f[457] && !f[373];
	assign leaf[13549] = !f[516] && f[544] && f[457] && f[373];
	assign leaf[13550] = f[516] && !f[601] && !f[660] && !f[295];
	assign leaf[13551] = f[516] && !f[601] && !f[660] && f[295];
	assign leaf[13552] = f[516] && !f[601] && f[660];
	assign leaf[13553] = f[516] && f[601] && !f[544];
	assign leaf[13554] = f[516] && f[601] && f[544] && !f[492];
	assign leaf[13555] = f[516] && f[601] && f[544] && f[492];
	
	// Tree 997, Classifier 7, Iteration: 99
	assign leaf[13556] = !f[396] && !f[376] && !f[288] && !f[261];
	assign leaf[13557] = !f[396] && !f[376] && !f[288] && f[261];
	assign leaf[13558] = !f[396] && !f[376] && f[288] && !f[290];
	assign leaf[13559] = !f[396] && !f[376] && f[288] && f[290];
	assign leaf[13560] = !f[396] && f[376] && !f[289] && !f[402];
	assign leaf[13561] = !f[396] && f[376] && !f[289] && f[402];
	assign leaf[13562] = !f[396] && f[376] && f[289] && !f[293];
	assign leaf[13563] = !f[396] && f[376] && f[289] && f[293];
	assign leaf[13564] = f[396] && !f[346] && !f[491];
	assign leaf[13565] = f[396] && !f[346] && f[491];
	assign leaf[13566] = f[396] && f[346];
	
	// Tree 998, Classifier 8, Iteration: 99
	assign leaf[13567] = !f[303] && !f[594] && !f[650] && !f[271];
	assign leaf[13568] = !f[303] && !f[594] && !f[650] && f[271];
	assign leaf[13569] = !f[303] && !f[594] && f[650] && !f[601];
	assign leaf[13570] = !f[303] && !f[594] && f[650] && f[601];
	assign leaf[13571] = !f[303] && f[594] && !f[463] && !f[465];
	assign leaf[13572] = !f[303] && f[594] && !f[463] && f[465];
	assign leaf[13573] = !f[303] && f[594] && f[463] && !f[487];
	assign leaf[13574] = !f[303] && f[594] && f[463] && f[487];
	assign leaf[13575] = f[303] && !f[649] && !f[682] && !f[207];
	assign leaf[13576] = f[303] && !f[649] && !f[682] && f[207];
	assign leaf[13577] = f[303] && !f[649] && f[682] && !f[595];
	assign leaf[13578] = f[303] && !f[649] && f[682] && f[595];
	assign leaf[13579] = f[303] && f[649];
	
	// Tree 999, Classifier 9, Iteration: 99
	assign leaf[13580] = !f[350] && !f[322] && !f[410] && !f[206];
	assign leaf[13581] = !f[350] && !f[322] && !f[410] && f[206];
	assign leaf[13582] = !f[350] && !f[322] && f[410] && !f[407];
	assign leaf[13583] = !f[350] && !f[322] && f[410] && f[407];
	assign leaf[13584] = !f[350] && f[322] && !f[266] && !f[352];
	assign leaf[13585] = !f[350] && f[322] && !f[266] && f[352];
	assign leaf[13586] = !f[350] && f[322] && f[266] && !f[238];
	assign leaf[13587] = !f[350] && f[322] && f[266] && f[238];
	assign leaf[13588] = f[350] && !f[324] && !f[430] && !f[204];
	assign leaf[13589] = f[350] && !f[324] && !f[430] && f[204];
	assign leaf[13590] = f[350] && !f[324] && f[430] && !f[211];
	assign leaf[13591] = f[350] && !f[324] && f[430] && f[211];
	assign leaf[13592] = f[350] && f[324] && !f[237] && !f[180];
	assign leaf[13593] = f[350] && f[324] && !f[237] && f[180];
	assign leaf[13594] = f[350] && f[324] && f[237] && !f[180];
	assign leaf[13595] = f[350] && f[324] && f[237] && f[180];
	
endmodule