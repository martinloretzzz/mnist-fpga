`timescale 1ns / 1ps

module leaf_counter_0(input logic [0:1411] l, output logic [7:0] val [0:12]);
	assign val[0] = l[0] + l[6] + l[12] + l[20] + l[24] + l[25] + l[27] + l[35] + l[39] + l[40] + l[42] + l[54] + l[67] + l[69] + l[73] + l[81] + l[85] + l[101] + l[106] + l[112] + l[116] + l[129] + l[132] + l[147] + l[151] + l[163] + l[166] + l[172] + l[182] + l[194] + l[200] + l[246] + l[259] + l[262] + l[275] + l[289] + l[313] + l[333] + l[339] + l[357] + l[364] + l[371] + l[375] + l[379] + l[385] + l[391] + l[398] + l[401] + l[429] + l[434] + l[440] + l[442] + l[444] + l[462] + l[468] + l[481] + l[489] + l[490] + l[494] + l[500] + l[505] + l[506] + l[508] + l[510] + l[527] + l[547] + l[565] + l[570] + l[575] + l[583] + l[596] + l[597] + l[603] + l[605] + l[623] + l[627] + l[643] + l[651] + l[668] + l[683] + l[688] + l[709] + l[759] + l[761] + l[763] + l[769] + l[780] + l[819] + l[844] + l[856] + l[861] + l[887] + l[909] + l[982] + l[984] + l[1009] + l[1014] + l[1063] + l[1073] + l[1086] + l[1145] + l[1213] + l[1237]; // -0.25
	assign val[1] = l[3] + l[13] + l[14] + l[18] + l[21] + l[22] + l[26] + l[33] + l[41] + l[43] + l[45] + l[48] + l[50] + l[52] + l[55] + l[57] + l[59] + l[61] + l[64] + l[70] + l[71] + l[72] + l[75] + l[83] + l[86] + l[88] + l[89] + l[93] + l[98] + l[102] + l[104] + l[110] + l[113] + l[114] + l[117] + l[119] + l[120] + l[123] + l[124] + l[126] + l[130] + l[133] + l[137] + l[140] + l[143] + l[145] + l[150] + l[155] + l[160] + l[164] + l[168] + l[171] + l[174] + l[178] + l[179] + l[180] + l[186] + l[188] + l[190] + l[202] + l[205] + l[206] + l[210] + l[211] + l[213] + l[215] + l[219] + l[221] + l[223] + l[225] + l[226] + l[230] + l[234] + l[235] + l[237] + l[239] + l[241] + l[242] + l[249] + l[251] + l[253] + l[258] + l[263] + l[265] + l[269] + l[273] + l[277] + l[282] + l[283] + l[285] + l[290] + l[291] + l[293] + l[296] + l[297] + l[300] + l[302] + l[303] + l[305] + l[309] + l[315] + l[317] + l[321] + l[327] + l[331] + l[335] + l[338] + l[341] + l[343] + l[345] + l[347] + l[349] + l[359] + l[365] + l[367] + l[369] + l[372] + l[381] + l[383] + l[386] + l[388] + l[395] + l[403] + l[407] + l[409] + l[412] + l[415] + l[423] + l[431] + l[433] + l[435] + l[443] + l[446] + l[447] + l[450] + l[454] + l[458] + l[461] + l[463] + l[465] + l[471] + l[472] + l[491] + l[492] + l[497] + l[502] + l[504] + l[517] + l[520] + l[522] + l[524] + l[529] + l[532] + l[533] + l[549] + l[552] + l[553] + l[558] + l[563] + l[568] + l[572] + l[573] + l[577] + l[580] + l[582] + l[589] + l[593] + l[606] + l[610] + l[612] + l[614] + l[626] + l[630] + l[634] + l[644] + l[648] + l[652] + l[656] + l[661] + l[663] + l[667] + l[670] + l[671] + l[673] + l[680] + l[682] + l[692] + l[694] + l[695] + l[698] + l[700] + l[704] + l[707] + l[712] + l[717] + l[723] + l[725] + l[727] + l[729] + l[730] + l[734] + l[737] + l[744] + l[746] + l[750] + l[772] + l[781] + l[786] + l[794] + l[795] + l[799] + l[800] + l[802] + l[806] + l[812] + l[813] + l[822] + l[826] + l[828] + l[835] + l[846] + l[850] + l[855] + l[862] + l[865] + l[870] + l[873] + l[878] + l[884] + l[891] + l[894] + l[895] + l[897] + l[905] + l[913] + l[918] + l[921] + l[929] + l[932] + l[933] + l[936] + l[937] + l[940] + l[944] + l[953] + l[960] + l[964] + l[966] + l[972] + l[977] + l[978] + l[981] + l[993] + l[995] + l[1011] + l[1027] + l[1030] + l[1033] + l[1039] + l[1040] + l[1042] + l[1044] + l[1046] + l[1047] + l[1055] + l[1057] + l[1059] + l[1062] + l[1066] + l[1068] + l[1072] + l[1077] + l[1080] + l[1084] + l[1089] + l[1093] + l[1098] + l[1099] + l[1101] + l[1111] + l[1118] + l[1122] + l[1123] + l[1130] + l[1131] + l[1136] + l[1142] + l[1143] + l[1146] + l[1152] + l[1154] + l[1161] + l[1166] + l[1167] + l[1174] + l[1179] + l[1181] + l[1187] + l[1190] + l[1198] + l[1199] + l[1209] + l[1217] + l[1223] + l[1228] + l[1233] + l[1240] + l[1246] + l[1255] + l[1256] + l[1258] + l[1263] + l[1270] + l[1274] + l[1283] + l[1287] + l[1293] + l[1300] + l[1308] + l[1310] + l[1316] + l[1320] + l[1327] + l[1330] + l[1335] + l[1337] + l[1344] + l[1352] + l[1358] + l[1368] + l[1378] + l[1385] + l[1399] + l[1408]; // -0.125
	assign val[2] = l[7] + l[29] + l[36] + l[37] + l[66] + l[77] + l[80] + l[82] + l[95] + l[107] + l[135] + l[148] + l[157] + l[162] + l[167] + l[176] + l[183] + l[185] + l[196] + l[214] + l[231] + l[247] + l[276] + l[279] + l[287] + l[326] + l[329] + l[354] + l[361] + l[374] + l[384] + l[390] + l[399] + l[404] + l[406] + l[414] + l[418] + l[419] + l[457] + l[470] + l[475] + l[476] + l[480] + l[487] + l[488] + l[499] + l[511] + l[513] + l[518] + l[525] + l[536] + l[538] + l[539] + l[541] + l[546] + l[569] + l[576] + l[585] + l[591] + l[595] + l[607] + l[615] + l[617] + l[625] + l[632] + l[639] + l[647] + l[650] + l[654] + l[659] + l[669] + l[675] + l[684] + l[686] + l[690] + l[710] + l[713] + l[715] + l[718] + l[719] + l[740] + l[742] + l[762] + l[767] + l[775] + l[784] + l[788] + l[791] + l[805] + l[809] + l[816] + l[820] + l[833] + l[836] + l[842] + l[860] + l[866] + l[871] + l[885] + l[900] + l[901] + l[906] + l[908] + l[914] + l[924] + l[945] + l[948] + l[949] + l[955] + l[958] + l[969] + l[998] + l[1000] + l[1005] + l[1007] + l[1010] + l[1019] + l[1028] + l[1050] + l[1054] + l[1060] + l[1075] + l[1083] + l[1096] + l[1106] + l[1113] + l[1133] + l[1139] + l[1141] + l[1155] + l[1156] + l[1163] + l[1172] + l[1188] + l[1191] + l[1203] + l[1206] + l[1211] + l[1212] + l[1214] + l[1227] + l[1229] + l[1232] + l[1238] + l[1251] + l[1254] + l[1260] + l[1267] + l[1277] + l[1282] + l[1289] + l[1298] + l[1305] + l[1318] + l[1333] + l[1340] + l[1346] + l[1353] + l[1359] + l[1362] + l[1366] + l[1369] + l[1375] + l[1379] + l[1382] + l[1387] + l[1392] + l[1393] + l[1396] + l[1404]; // -0.0625
	assign val[3] = l[28] + l[90] + l[121] + l[134] + l[138] + l[152] + l[153] + l[227] + l[245] + l[255] + l[272] + l[292] + l[312] + l[334] + l[351] + l[358] + l[366] + l[397] + l[484] + l[501] + l[548] + l[555] + l[566] + l[588] + l[600] + l[636] + l[674] + l[677] + l[687] + l[696] + l[722] + l[728] + l[749] + l[774] + l[779] + l[807] + l[810] + l[814] + l[817] + l[830] + l[841] + l[847] + l[854] + l[858] + l[876] + l[882] + l[888] + l[898] + l[930] + l[951] + l[967] + l[979] + l[985] + l[986] + l[990] + l[1023] + l[1024] + l[1032] + l[1036] + l[1041] + l[1064] + l[1067] + l[1091] + l[1108] + l[1121] + l[1149] + l[1151] + l[1153] + l[1178] + l[1194] + l[1220] + l[1235] + l[1243] + l[1248] + l[1264] + l[1284] + l[1311] + l[1314] + l[1315] + l[1321] + l[1322] + l[1326] + l[1332] + l[1355] + l[1361] + l[1365] + l[1390] + l[1394] + l[1406]; // -0.03125
	assign val[4] = l[74] + l[87] + l[118] + l[192] + l[217] + l[243] + l[267] + l[314] + l[323] + l[394] + l[428] + l[452] + l[469] + l[495] + l[528] + l[609] + l[619] + l[624] + l[629] + l[635] + l[837] + l[874] + l[879] + l[910] + l[927] + l[963] + l[974] + l[1021] + l[1034] + l[1094] + l[1110] + l[1115] + l[1127] + l[1175] + l[1202] + l[1215] + l[1231] + l[1242] + l[1329] + l[1338] + l[1345] + l[1400]; // -0.015625
	assign val[5] = l[56] + l[58] + l[199] + l[266] + l[274] + l[356] + l[377] + l[411] + l[455] + l[464] + l[485] + l[571] + l[581] + l[657] + l[662] + l[697] + l[783] + l[793] + l[808] + l[815] + l[823] + l[863] + l[883] + l[904] + l[912] + l[976] + l[980] + l[996] + l[1013] + l[1052] + l[1056] + l[1097] + l[1119] + l[1129] + l[1150] + l[1200] + l[1207] + l[1224] + l[1245] + l[1257] + l[1276] + l[1281] + l[1291] + l[1294] + l[1317] + l[1328] + l[1342] + l[1349] + l[1367] + l[1370] + l[1381] + l[1409]; // 0.015625
	assign val[6] = l[131] + l[220] + l[260] + l[284] + l[295] + l[318] + l[332] + l[350] + l[362] + l[368] + l[416] + l[421] + l[424] + l[445] + l[477] + l[493] + l[498] + l[507] + l[509] + l[514] + l[521] + l[534] + l[537] + l[557] + l[590] + l[618] + l[640] + l[664] + l[679] + l[691] + l[720] + l[726] + l[738] + l[741] + l[743] + l[747] + l[770] + l[796] + l[818] + l[821] + l[840] + l[872] + l[892] + l[902] + l[939] + l[942] + l[959] + l[973] + l[983] + l[988] + l[997] + l[1049] + l[1053] + l[1058] + l[1061] + l[1079] + l[1085] + l[1090] + l[1105] + l[1117] + l[1137] + l[1140] + l[1164] + l[1168] + l[1193] + l[1196] + l[1204] + l[1210] + l[1230] + l[1259] + l[1262] + l[1266] + l[1271] + l[1272] + l[1295] + l[1301] + l[1304] + l[1324] + l[1334] + l[1341] + l[1377] + l[1391] + l[1397] + l[1405] + l[1410]; // 0.03125
	assign val[7] = l[108] + l[111] + l[141] + l[159] + l[173] + l[208] + l[212] + l[224] + l[250] + l[257] + l[270] + l[286] + l[316] + l[322] + l[337] + l[340] + l[342] + l[363] + l[380] + l[396] + l[410] + l[430] + l[449] + l[456] + l[459] + l[474] + l[483] + l[503] + l[526] + l[530] + l[531] + l[542] + l[545] + l[554] + l[567] + l[578] + l[579] + l[604] + l[611] + l[620] + l[637] + l[660] + l[672] + l[685] + l[693] + l[699] + l[711] + l[721] + l[731] + l[732] + l[735] + l[736] + l[745] + l[751] + l[764] + l[768] + l[773] + l[776] + l[782] + l[798] + l[803] + l[804] + l[811] + l[824] + l[827] + l[831] + l[832] + l[834] + l[839] + l[853] + l[864] + l[886] + l[893] + l[907] + l[915] + l[916] + l[925] + l[934] + l[935] + l[950] + l[954] + l[962] + l[968] + l[987] + l[992] + l[999] + l[1002] + l[1004] + l[1006] + l[1022] + l[1031] + l[1035] + l[1038] + l[1043] + l[1045] + l[1048] + l[1071] + l[1076] + l[1081] + l[1092] + l[1095] + l[1102] + l[1109] + l[1112] + l[1128] + l[1134] + l[1157] + l[1159] + l[1162] + l[1165] + l[1169] + l[1173] + l[1176] + l[1177] + l[1180] + l[1182] + l[1185] + l[1192] + l[1205] + l[1208] + l[1218] + l[1219] + l[1234] + l[1241] + l[1244] + l[1247] + l[1252] + l[1265] + l[1278] + l[1288] + l[1290] + l[1299] + l[1306] + l[1312] + l[1313] + l[1319] + l[1331] + l[1339] + l[1347] + l[1351] + l[1354] + l[1356] + l[1360] + l[1376] + l[1389] + l[1395] + l[1407]; // 0.0625
	assign val[8] = l[4] + l[16] + l[31] + l[34] + l[46] + l[49] + l[51] + l[53] + l[62] + l[68] + l[94] + l[97] + l[100] + l[103] + l[122] + l[125] + l[127] + l[139] + l[144] + l[146] + l[156] + l[161] + l[169] + l[170] + l[177] + l[189] + l[191] + l[193] + l[195] + l[197] + l[201] + l[204] + l[207] + l[209] + l[218] + l[233] + l[236] + l[240] + l[248] + l[256] + l[261] + l[264] + l[268] + l[280] + l[281] + l[288] + l[298] + l[299] + l[301] + l[304] + l[308] + l[310] + l[311] + l[320] + l[328] + l[330] + l[344] + l[348] + l[352] + l[353] + l[360] + l[373] + l[378] + l[382] + l[387] + l[389] + l[393] + l[400] + l[405] + l[413] + l[417] + l[420] + l[422] + l[426] + l[427] + l[432] + l[439] + l[453] + l[460] + l[466] + l[473] + l[479] + l[486] + l[496] + l[519] + l[523] + l[535] + l[551] + l[556] + l[560] + l[562] + l[574] + l[586] + l[587] + l[592] + l[594] + l[599] + l[602] + l[613] + l[616] + l[621] + l[633] + l[638] + l[642] + l[645] + l[646] + l[649] + l[653] + l[655] + l[658] + l[665] + l[666] + l[676] + l[678] + l[706] + l[708] + l[716] + l[739] + l[748] + l[753] + l[756] + l[758] + l[766] + l[785] + l[787] + l[792] + l[843] + l[849] + l[859] + l[867] + l[868] + l[875] + l[880] + l[881] + l[890] + l[896] + l[899] + l[903] + l[911] + l[922] + l[926] + l[931] + l[946] + l[947] + l[952] + l[970] + l[975] + l[989] + l[1008] + l[1016] + l[1020] + l[1025] + l[1029] + l[1037] + l[1051] + l[1065] + l[1070] + l[1078] + l[1082] + l[1088] + l[1104] + l[1107] + l[1114] + l[1116] + l[1125] + l[1138] + l[1148] + l[1158] + l[1170] + l[1184] + l[1195] + l[1201] + l[1216] + l[1222] + l[1226] + l[1249] + l[1253] + l[1261] + l[1269] + l[1275] + l[1279] + l[1285] + l[1292] + l[1296] + l[1302] + l[1323] + l[1325] + l[1343] + l[1350] + l[1364] + l[1372] + l[1373] + l[1383] + l[1398] + l[1401] + l[1403] + l[1411]; // 0.125
	assign val[9] = l[8] + l[11] + l[19] + l[23] + l[38] + l[44] + l[47] + l[60] + l[63] + l[65] + l[76] + l[78] + l[79] + l[84] + l[96] + l[99] + l[109] + l[115] + l[128] + l[136] + l[142] + l[158] + l[181] + l[184] + l[198] + l[216] + l[228] + l[232] + l[244] + l[252] + l[271] + l[294] + l[324] + l[325] + l[355] + l[437] + l[451] + l[478] + l[512] + l[516] + l[540] + l[543] + l[608] + l[628] + l[641] + l[689] + l[702] + l[714] + l[733] + l[755] + l[777] + l[790] + l[797] + l[825] + l[838] + l[917] + l[941] + l[956] + l[1001] + l[1120]; // 0.25
	assign val[10] = l[15] + l[17] + l[30] + l[32] + l[91] + l[105] + l[154]; // 0.5
	assign val[11] = l[2] + l[5] + l[9]; // 1.0
	assign val[12] = l[10]; // 2.0
endmodule

module leaf_counter_1(input logic [0:1154] l, output logic [7:0] val [0:12]);
	assign val[0] = l[0] + l[2] + l[4] + l[5] + l[7] + l[15] + l[21] + l[23] + l[27] + l[34] + l[36] + l[37] + l[41] + l[45] + l[46] + l[50] + l[54] + l[57] + l[61] + l[63] + l[65] + l[71] + l[80] + l[82] + l[84] + l[85] + l[92] + l[94] + l[95] + l[101] + l[107] + l[110] + l[111] + l[118] + l[127] + l[128] + l[131] + l[134] + l[136] + l[142] + l[148] + l[152] + l[153] + l[162] + l[164] + l[168] + l[172] + l[173] + l[182] + l[187] + l[188] + l[192] + l[198] + l[199] + l[201] + l[203] + l[205] + l[210] + l[219] + l[220] + l[224] + l[228] + l[230] + l[232] + l[233] + l[243] + l[244] + l[254] + l[257] + l[258] + l[266] + l[270] + l[272] + l[278] + l[279] + l[282] + l[284] + l[285] + l[288] + l[290] + l[296] + l[300] + l[304] + l[307] + l[314] + l[316] + l[317] + l[319] + l[322] + l[327] + l[328] + l[333] + l[337] + l[341] + l[342] + l[352] + l[357] + l[359] + l[360] + l[368] + l[369] + l[376] + l[377] + l[382] + l[389] + l[392] + l[397] + l[398] + l[400] + l[402] + l[405] + l[407] + l[408] + l[412] + l[418] + l[420] + l[421] + l[433] + l[437] + l[442] + l[447] + l[449] + l[450] + l[459] + l[460] + l[463] + l[464] + l[468] + l[476] + l[478] + l[484] + l[488] + l[491] + l[493] + l[496] + l[501] + l[502] + l[507] + l[513] + l[519] + l[523] + l[526] + l[528] + l[534] + l[536] + l[539] + l[546] + l[553] + l[556] + l[557] + l[559] + l[560] + l[572] + l[578] + l[584] + l[590] + l[596] + l[599] + l[602] + l[603] + l[612] + l[621] + l[623] + l[632] + l[636] + l[639] + l[643] + l[645] + l[653] + l[665] + l[673] + l[676] + l[679] + l[683] + l[692] + l[694] + l[697] + l[700] + l[705] + l[707] + l[713] + l[716] + l[730] + l[737] + l[739] + l[747] + l[749] + l[754] + l[766] + l[779] + l[797] + l[800] + l[811] + l[823] + l[825] + l[839] + l[844] + l[853] + l[859] + l[866] + l[872] + l[888] + l[890] + l[891] + l[894] + l[907] + l[932] + l[947] + l[964] + l[965] + l[974] + l[984] + l[989] + l[991] + l[995] + l[1013] + l[1021] + l[1038] + l[1040] + l[1057] + l[1085] + l[1100] + l[1110] + l[1118] + l[1130] + l[1140] + l[1141]; // -0.25
	assign val[1] = l[1] + l[6] + l[10] + l[14] + l[16] + l[18] + l[24] + l[25] + l[30] + l[31] + l[33] + l[38] + l[39] + l[42] + l[44] + l[48] + l[49] + l[52] + l[55] + l[58] + l[60] + l[68] + l[69] + l[73] + l[74] + l[77] + l[78] + l[83] + l[88] + l[89] + l[91] + l[96] + l[98] + l[100] + l[104] + l[108] + l[113] + l[115] + l[116] + l[119] + l[120] + l[122] + l[126] + l[130] + l[133] + l[138] + l[140] + l[141] + l[143] + l[145] + l[154] + l[156] + l[157] + l[159] + l[166] + l[167] + l[174] + l[175] + l[177] + l[179] + l[191] + l[193] + l[196] + l[204] + l[208] + l[212] + l[215] + l[217] + l[221] + l[223] + l[226] + l[229] + l[235] + l[246] + l[247] + l[248] + l[250] + l[253] + l[259] + l[267] + l[268] + l[271] + l[273] + l[275] + l[281] + l[292] + l[293] + l[302] + l[305] + l[309] + l[311] + l[325] + l[331] + l[334] + l[339] + l[344] + l[347] + l[348] + l[350] + l[354] + l[356] + l[363] + l[367] + l[371] + l[378] + l[381] + l[383] + l[386] + l[391] + l[395] + l[415] + l[424] + l[428] + l[431] + l[435] + l[439] + l[440] + l[448] + l[451] + l[455] + l[462] + l[467] + l[469] + l[471] + l[481] + l[492] + l[495] + l[503] + l[505] + l[509] + l[515] + l[517] + l[520] + l[524] + l[527] + l[529] + l[537] + l[544] + l[570] + l[573] + l[580] + l[587] + l[593] + l[604] + l[609] + l[617] + l[618] + l[627] + l[629] + l[631] + l[634] + l[647] + l[651] + l[654] + l[656] + l[658] + l[661] + l[662] + l[666] + l[671] + l[674] + l[684] + l[688] + l[690] + l[693] + l[695] + l[703] + l[710] + l[718] + l[723] + l[724] + l[726] + l[727] + l[732] + l[740] + l[744] + l[746] + l[748] + l[750] + l[758] + l[762] + l[763] + l[765] + l[769] + l[772] + l[777] + l[785] + l[787] + l[793] + l[794] + l[799] + l[803] + l[817] + l[820] + l[822] + l[830] + l[834] + l[836] + l[838] + l[841] + l[851] + l[856] + l[863] + l[865] + l[868] + l[870] + l[873] + l[874] + l[882] + l[904] + l[905] + l[909] + l[910] + l[913] + l[916] + l[924] + l[925] + l[928] + l[929] + l[931] + l[934] + l[936] + l[937] + l[940] + l[950] + l[956] + l[957] + l[959] + l[969] + l[972] + l[980] + l[983] + l[993] + l[996] + l[1001] + l[1004] + l[1007] + l[1009] + l[1011] + l[1014] + l[1016] + l[1025] + l[1032] + l[1034] + l[1044] + l[1046] + l[1049] + l[1055] + l[1060] + l[1062] + l[1066] + l[1070] + l[1073] + l[1077] + l[1086] + l[1089] + l[1091] + l[1094] + l[1102] + l[1104] + l[1106] + l[1114] + l[1122] + l[1125] + l[1132] + l[1137] + l[1143] + l[1151]; // -0.125
	assign val[2] = l[8] + l[20] + l[28] + l[29] + l[35] + l[43] + l[53] + l[64] + l[66] + l[75] + l[81] + l[86] + l[102] + l[112] + l[121] + l[161] + l[183] + l[184] + l[189] + l[206] + l[211] + l[231] + l[238] + l[274] + l[287] + l[298] + l[303] + l[308] + l[330] + l[332] + l[345] + l[353] + l[364] + l[370] + l[374] + l[375] + l[387] + l[393] + l[401] + l[403] + l[411] + l[422] + l[436] + l[473] + l[489] + l[499] + l[512] + l[543] + l[548] + l[561] + l[563] + l[566] + l[569] + l[577] + l[585] + l[589] + l[591] + l[598] + l[607] + l[611] + l[613] + l[625] + l[642] + l[644] + l[646] + l[664] + l[672] + l[678] + l[681] + l[687] + l[712] + l[715] + l[720] + l[729] + l[735] + l[742] + l[751] + l[759] + l[782] + l[784] + l[796] + l[807] + l[810] + l[816] + l[826] + l[845] + l[850] + l[880] + l[892] + l[893] + l[901] + l[914] + l[918] + l[920] + l[941] + l[951] + l[953] + l[1018] + l[1024] + l[1028] + l[1029] + l[1039] + l[1051] + l[1058] + l[1072] + l[1081] + l[1082] + l[1084] + l[1093] + l[1107] + l[1112] + l[1119] + l[1139]; // -0.0625
	assign val[3] = l[109] + l[129] + l[186] + l[207] + l[213] + l[236] + l[313] + l[318] + l[321] + l[329] + l[336] + l[361] + l[458] + l[465] + l[475] + l[506] + l[510] + l[531] + l[535] + l[558] + l[581] + l[624] + l[704] + l[731] + l[756] + l[774] + l[778] + l[788] + l[808] + l[814] + l[842] + l[848] + l[854] + l[855] + l[877] + l[879] + l[883] + l[887] + l[900] + l[912] + l[935] + l[944] + l[945] + l[960] + l[962] + l[963] + l[966] + l[975] + l[985] + l[988] + l[990] + l[1010] + l[1022] + l[1037] + l[1042] + l[1043] + l[1048] + l[1052] + l[1056] + l[1064] + l[1080] + l[1099] + l[1113] + l[1121] + l[1127] + l[1129] + l[1142] + l[1148] + l[1152]; // -0.03125
	assign val[4] = l[22] + l[67] + l[149] + l[200] + l[245] + l[264] + l[324] + l[340] + l[417] + l[427] + l[444] + l[470] + l[533] + l[635] + l[659] + l[706] + l[767] + l[773] + l[818] + l[829] + l[933] + l[948] + l[978] + l[1036] + l[1074] + l[1115]; // -0.015625
	assign val[5] = l[79] + l[137] + l[222] + l[242] + l[294] + l[301] + l[438] + l[454] + l[461] + l[474] + l[582] + l[594] + l[622] + l[691] + l[728] + l[753] + l[757] + l[864] + l[871] + l[895] + l[952] + l[992] + l[994] + l[1071] + l[1103] + l[1117] + l[1144]; // 0.015625
	assign val[6] = l[62] + l[70] + l[72] + l[117] + l[146] + l[180] + l[225] + l[277] + l[286] + l[315] + l[373] + l[423] + l[429] + l[432] + l[445] + l[452] + l[453] + l[479] + l[498] + l[522] + l[547] + l[554] + l[568] + l[605] + l[641] + l[667] + l[677] + l[711] + l[722] + l[760] + l[764] + l[768] + l[775] + l[791] + l[812] + l[824] + l[828] + l[835] + l[840] + l[849] + l[889] + l[967] + l[976] + l[979] + l[1003] + l[1012] + l[1023] + l[1054] + l[1088] + l[1095] + l[1128] + l[1133] + l[1147] + l[1149]; // 0.03125
	assign val[7] = l[40] + l[90] + l[147] + l[151] + l[163] + l[185] + l[195] + l[197] + l[202] + l[218] + l[234] + l[252] + l[255] + l[256] + l[283] + l[295] + l[312] + l[323] + l[335] + l[355] + l[362] + l[379] + l[384] + l[385] + l[394] + l[396] + l[399] + l[404] + l[410] + l[414] + l[416] + l[426] + l[434] + l[441] + l[446] + l[482] + l[494] + l[500] + l[504] + l[516] + l[521] + l[530] + l[532] + l[540] + l[574] + l[586] + l[620] + l[626] + l[633] + l[640] + l[648] + l[650] + l[657] + l[669] + l[675] + l[686] + l[696] + l[699] + l[701] + l[702] + l[717] + l[725] + l[736] + l[741] + l[745] + l[770] + l[792] + l[798] + l[819] + l[821] + l[832] + l[852] + l[861] + l[867] + l[869] + l[899] + l[902] + l[927] + l[943] + l[961] + l[981] + l[982] + l[1002] + l[1008] + l[1017] + l[1033] + l[1035] + l[1041] + l[1047] + l[1053] + l[1061] + l[1083] + l[1090] + l[1105] + l[1111] + l[1126] + l[1136] + l[1153]; // 0.0625
	assign val[8] = l[26] + l[47] + l[56] + l[97] + l[99] + l[103] + l[105] + l[114] + l[123] + l[125] + l[132] + l[135] + l[139] + l[144] + l[150] + l[160] + l[171] + l[181] + l[216] + l[227] + l[240] + l[262] + l[265] + l[269] + l[280] + l[291] + l[299] + l[306] + l[346] + l[349] + l[358] + l[372] + l[380] + l[388] + l[390] + l[406] + l[457] + l[466] + l[487] + l[511] + l[514] + l[525] + l[538] + l[545] + l[562] + l[567] + l[579] + l[592] + l[595] + l[614] + l[630] + l[637] + l[655] + l[680] + l[682] + l[689] + l[709] + l[733] + l[734] + l[738] + l[743] + l[752] + l[755] + l[776] + l[781] + l[783] + l[795] + l[805] + l[809] + l[815] + l[843] + l[847] + l[857] + l[862] + l[875] + l[876] + l[878] + l[885] + l[896] + l[898] + l[903] + l[915] + l[930] + l[938] + l[939] + l[942] + l[946] + l[949] + l[954] + l[955] + l[968] + l[973] + l[977] + l[986] + l[987] + l[998] + l[1006] + l[1015] + l[1019] + l[1031] + l[1059] + l[1063] + l[1067] + l[1068] + l[1079] + l[1087] + l[1092] + l[1097] + l[1101] + l[1108] + l[1116] + l[1120] + l[1123] + l[1131] + l[1134] + l[1145] + l[1154]; // 0.125
	assign val[9] = l[3] + l[13] + l[51] + l[59] + l[76] + l[93] + l[106] + l[155] + l[176] + l[178] + l[190] + l[209] + l[237] + l[251] + l[263] + l[276] + l[310] + l[320] + l[351] + l[365] + l[409] + l[425] + l[472] + l[483] + l[541] + l[549] + l[551] + l[565] + l[575] + l[583] + l[588] + l[606] + l[610] + l[615] + l[619] + l[628] + l[638] + l[649] + l[663] + l[670] + l[685] + l[698] + l[719] + l[721] + l[761] + l[771] + l[780] + l[789] + l[813] + l[827] + l[833] + l[884] + l[919] + l[921] + l[971] + l[1000] + l[1027] + l[1050] + l[1075] + l[1098] + l[1150]; // 0.25
	assign val[10] = l[19] + l[32] + l[87] + l[214] + l[239] + l[297] + l[480] + l[485] + l[550] + l[564] + l[576] + l[790] + l[897]; // 0.5
	assign val[11] = l[9] + l[11]; // 1.0
	assign val[12] = 0; // 2.0
endmodule

module leaf_counter_2(input logic [0:1374] l, output logic [7:0] val [0:12]);
	assign val[0] = l[12] + l[38] + l[51] + l[61] + l[71] + l[98] + l[109] + l[139] + l[145] + l[184] + l[185] + l[232] + l[238] + l[257] + l[262] + l[263] + l[281] + l[298] + l[305] + l[323] + l[329] + l[342] + l[350] + l[371] + l[394] + l[409] + l[411] + l[423] + l[450] + l[467] + l[469] + l[473] + l[484] + l[490] + l[501] + l[505] + l[509] + l[510] + l[511] + l[517] + l[522] + l[535] + l[551] + l[575] + l[591] + l[596] + l[606] + l[610] + l[618] + l[621] + l[654] + l[656] + l[667] + l[678] + l[702] + l[706] + l[708] + l[725] + l[740] + l[742] + l[757] + l[804] + l[808] + l[839] + l[844] + l[850] + l[867] + l[882] + l[896] + l[963] + l[965] + l[978] + l[994] + l[1031] + l[1033] + l[1042] + l[1055] + l[1071] + l[1073] + l[1080] + l[1084] + l[1089] + l[1103] + l[1116] + l[1145] + l[1168] + l[1189] + l[1235] + l[1248] + l[1322]; // -0.25
	assign val[1] = l[0] + l[6] + l[16] + l[17] + l[21] + l[22] + l[27] + l[28] + l[31] + l[32] + l[35] + l[40] + l[43] + l[48] + l[53] + l[54] + l[56] + l[67] + l[72] + l[75] + l[79] + l[84] + l[86] + l[90] + l[94] + l[95] + l[100] + l[103] + l[113] + l[118] + l[119] + l[121] + l[126] + l[129] + l[131] + l[140] + l[146] + l[149] + l[150] + l[152] + l[154] + l[157] + l[162] + l[164] + l[169] + l[171] + l[174] + l[179] + l[180] + l[188] + l[189] + l[195] + l[202] + l[208] + l[209] + l[212] + l[213] + l[218] + l[219] + l[225] + l[228] + l[229] + l[233] + l[239] + l[244] + l[246] + l[247] + l[249] + l[258] + l[265] + l[269] + l[271] + l[280] + l[287] + l[294] + l[295] + l[301] + l[307] + l[310] + l[313] + l[317] + l[325] + l[334] + l[340] + l[348] + l[358] + l[361] + l[365] + l[367] + l[368] + l[375] + l[377] + l[380] + l[383] + l[389] + l[399] + l[400] + l[417] + l[421] + l[424] + l[430] + l[432] + l[434] + l[440] + l[443] + l[444] + l[446] + l[466] + l[475] + l[482] + l[498] + l[502] + l[527] + l[529] + l[544] + l[548] + l[550] + l[555] + l[559] + l[569] + l[577] + l[578] + l[580] + l[585] + l[589] + l[602] + l[616] + l[631] + l[634] + l[636] + l[638] + l[643] + l[646] + l[649] + l[665] + l[669] + l[683] + l[686] + l[695] + l[697] + l[701] + l[720] + l[724] + l[727] + l[736] + l[745] + l[751] + l[753] + l[760] + l[762] + l[766] + l[779] + l[780] + l[782] + l[784] + l[788] + l[792] + l[795] + l[797] + l[798] + l[803] + l[811] + l[816] + l[818] + l[820] + l[824] + l[833] + l[837] + l[843] + l[857] + l[863] + l[869] + l[870] + l[875] + l[889] + l[891] + l[901] + l[904] + l[905] + l[908] + l[911] + l[920] + l[924] + l[926] + l[928] + l[931] + l[939] + l[941] + l[944] + l[946] + l[948] + l[955] + l[957] + l[960] + l[971] + l[979] + l[986] + l[1003] + l[1005] + l[1006] + l[1016] + l[1021] + l[1022] + l[1038] + l[1044] + l[1045] + l[1059] + l[1067] + l[1070] + l[1075] + l[1079] + l[1087] + l[1091] + l[1097] + l[1106] + l[1109] + l[1120] + l[1122] + l[1123] + l[1128] + l[1134] + l[1144] + l[1150] + l[1151] + l[1161] + l[1164] + l[1166] + l[1172] + l[1178] + l[1179] + l[1181] + l[1182] + l[1191] + l[1200] + l[1205] + l[1206] + l[1212] + l[1218] + l[1222] + l[1227] + l[1232] + l[1237] + l[1242] + l[1245] + l[1251] + l[1262] + l[1270] + l[1278] + l[1284] + l[1286] + l[1300] + l[1301] + l[1307] + l[1314] + l[1315] + l[1330] + l[1333] + l[1339] + l[1349] + l[1351] + l[1353] + l[1355] + l[1357] + l[1358] + l[1363] + l[1369]; // -0.125
	assign val[2] = l[15] + l[18] + l[37] + l[46] + l[63] + l[73] + l[82] + l[102] + l[106] + l[115] + l[134] + l[137] + l[153] + l[158] + l[161] + l[166] + l[177] + l[196] + l[199] + l[204] + l[221] + l[243] + l[251] + l[254] + l[255] + l[273] + l[283] + l[289] + l[327] + l[330] + l[331] + l[337] + l[343] + l[344] + l[352] + l[354] + l[357] + l[370] + l[378] + l[390] + l[396] + l[404] + l[410] + l[413] + l[414] + l[422] + l[454] + l[457] + l[459] + l[462] + l[472] + l[479] + l[489] + l[491] + l[493] + l[504] + l[514] + l[515] + l[523] + l[530] + l[531] + l[536] + l[560] + l[563] + l[567] + l[571] + l[573] + l[583] + l[587] + l[620] + l[622] + l[625] + l[628] + l[650] + l[661] + l[663] + l[668] + l[676] + l[682] + l[689] + l[709] + l[715] + l[723] + l[731] + l[735] + l[747] + l[756] + l[768] + l[771] + l[815] + l[823] + l[838] + l[845] + l[846] + l[851] + l[852] + l[858] + l[861] + l[876] + l[879] + l[880] + l[890] + l[893] + l[897] + l[900] + l[907] + l[913] + l[929] + l[935] + l[949] + l[969] + l[976] + l[983] + l[993] + l[997] + l[998] + l[1001] + l[1010] + l[1013] + l[1014] + l[1020] + l[1026] + l[1032] + l[1034] + l[1040] + l[1043] + l[1077] + l[1082] + l[1085] + l[1095] + l[1115] + l[1130] + l[1153] + l[1154] + l[1159] + l[1184] + l[1187] + l[1193] + l[1213] + l[1220] + l[1225] + l[1234] + l[1254] + l[1257] + l[1258] + l[1264] + l[1276] + l[1281] + l[1283] + l[1289] + l[1309] + l[1312] + l[1319] + l[1321] + l[1325] + l[1327] + l[1338] + l[1366] + l[1367] + l[1372]; // -0.0625
	assign val[3] = l[39] + l[85] + l[87] + l[91] + l[117] + l[170] + l[186] + l[191] + l[226] + l[242] + l[264] + l[278] + l[282] + l[288] + l[297] + l[315] + l[381] + l[387] + l[407] + l[436] + l[452] + l[474] + l[487] + l[495] + l[507] + l[533] + l[542] + l[584] + l[605] + l[609] + l[611] + l[648] + l[677] + l[680] + l[694] + l[729] + l[741] + l[744] + l[754] + l[774] + l[787] + l[791] + l[800] + l[809] + l[812] + l[840] + l[854] + l[856] + l[862] + l[883] + l[884] + l[895] + l[918] + l[932] + l[945] + l[974] + l[981] + l[991] + l[1023] + l[1049] + l[1051] + l[1064] + l[1092] + l[1101] + l[1104] + l[1118] + l[1131] + l[1137] + l[1158] + l[1174] + l[1197] + l[1199] + l[1207] + l[1217] + l[1229] + l[1230] + l[1240] + l[1261] + l[1279] + l[1291] + l[1294] + l[1304] + l[1305] + l[1318] + l[1329] + l[1336] + l[1344] + l[1347] + l[1348]; // -0.03125
	assign val[4] = l[57] + l[80] + l[173] + l[306] + l[435] + l[439] + l[477] + l[486] + l[526] + l[552] + l[592] + l[599] + l[619] + l[640] + l[660] + l[671] + l[739] + l[773] + l[777] + l[781] + l[794] + l[806] + l[807] + l[830] + l[887] + l[910] + l[914] + l[933] + l[987] + l[995] + l[1056] + l[1060] + l[1061] + l[1074] + l[1090] + l[1110] + l[1133] + l[1185] + l[1216] + l[1241] + l[1268] + l[1334] + l[1340]; // -0.015625
	assign val[5] = l[78] + l[107] + l[151] + l[215] + l[237] + l[261] + l[272] + l[318] + l[322] + l[341] + l[416] + l[418] + l[441] + l[516] + l[518] + l[538] + l[556] + l[574] + l[612] + l[655] + l[692] + l[696] + l[728] + l[737] + l[750] + l[752] + l[834] + l[853] + l[865] + l[868] + l[871] + l[902] + l[951] + l[953] + l[958] + l[972] + l[975] + l[980] + l[1019] + l[1039] + l[1052] + l[1057] + l[1081] + l[1088] + l[1096] + l[1102] + l[1108] + l[1112] + l[1114] + l[1124] + l[1125] + l[1192] + l[1196] + l[1224] + l[1228] + l[1296] + l[1326] + l[1370]; // 0.015625
	assign val[6] = l[5] + l[125] + l[143] + l[205] + l[224] + l[235] + l[285] + l[304] + l[319] + l[366] + l[369] + l[425] + l[442] + l[449] + l[456] + l[465] + l[468] + l[506] + l[521] + l[540] + l[541] + l[543] + l[566] + l[588] + l[590] + l[632] + l[644] + l[693] + l[698] + l[730] + l[764] + l[767] + l[770] + l[805] + l[826] + l[866] + l[898] + l[906] + l[916] + l[930] + l[943] + l[964] + l[967] + l[990] + l[1002] + l[1004] + l[1007] + l[1008] + l[1012] + l[1078] + l[1098] + l[1100] + l[1121] + l[1155] + l[1160] + l[1183] + l[1198] + l[1201] + l[1208] + l[1210] + l[1211] + l[1239] + l[1247] + l[1250] + l[1263] + l[1274] + l[1280] + l[1303] + l[1320] + l[1337] + l[1352] + l[1371]; // 0.03125
	assign val[7] = l[3] + l[41] + l[62] + l[111] + l[181] + l[198] + l[207] + l[220] + l[222] + l[240] + l[250] + l[260] + l[314] + l[338] + l[346] + l[349] + l[351] + l[359] + l[360] + l[376] + l[388] + l[391] + l[392] + l[395] + l[420] + l[445] + l[451] + l[453] + l[458] + l[463] + l[480] + l[481] + l[496] + l[503] + l[512] + l[513] + l[524] + l[525] + l[576] + l[579] + l[586] + l[600] + l[604] + l[615] + l[617] + l[623] + l[624] + l[652] + l[659] + l[664] + l[699] + l[703] + l[710] + l[714] + l[743] + l[746] + l[761] + l[772] + l[775] + l[783] + l[790] + l[793] + l[799] + l[801] + l[802] + l[810] + l[814] + l[821] + l[822] + l[825] + l[848] + l[860] + l[864] + l[874] + l[877] + l[881] + l[899] + l[921] + l[922] + l[927] + l[934] + l[940] + l[947] + l[962] + l[985] + l[989] + l[992] + l[1000] + l[1011] + l[1018] + l[1027] + l[1028] + l[1036] + l[1046] + l[1047] + l[1068] + l[1069] + l[1093] + l[1094] + l[1107] + l[1140] + l[1148] + l[1149] + l[1152] + l[1156] + l[1162] + l[1169] + l[1186] + l[1188] + l[1194] + l[1215] + l[1223] + l[1226] + l[1246] + l[1252] + l[1256] + l[1260] + l[1265] + l[1269] + l[1277] + l[1282] + l[1287] + l[1290] + l[1292] + l[1293] + l[1297] + l[1306] + l[1310] + l[1311] + l[1316] + l[1317] + l[1323] + l[1331] + l[1335] + l[1341] + l[1345] + l[1350] + l[1354] + l[1356] + l[1359] + l[1361] + l[1368]; // 0.0625
	assign val[8] = l[9] + l[13] + l[26] + l[29] + l[59] + l[65] + l[68] + l[96] + l[97] + l[99] + l[104] + l[128] + l[130] + l[156] + l[159] + l[160] + l[163] + l[167] + l[192] + l[217] + l[223] + l[227] + l[245] + l[248] + l[252] + l[253] + l[266] + l[268] + l[274] + l[279] + l[284] + l[291] + l[293] + l[300] + l[302] + l[303] + l[308] + l[316] + l[332] + l[336] + l[345] + l[347] + l[355] + l[363] + l[384] + l[393] + l[397] + l[398] + l[403] + l[405] + l[406] + l[408] + l[415] + l[419] + l[427] + l[433] + l[438] + l[447] + l[448] + l[455] + l[461] + l[471] + l[478] + l[483] + l[488] + l[494] + l[497] + l[500] + l[508] + l[532] + l[537] + l[547] + l[549] + l[554] + l[557] + l[561] + l[565] + l[570] + l[572] + l[581] + l[582] + l[595] + l[598] + l[607] + l[613] + l[626] + l[629] + l[630] + l[633] + l[637] + l[641] + l[647] + l[651] + l[658] + l[662] + l[672] + l[675] + l[679] + l[688] + l[690] + l[718] + l[722] + l[726] + l[733] + l[738] + l[749] + l[755] + l[758] + l[769] + l[776] + l[786] + l[796] + l[817] + l[819] + l[827] + l[831] + l[835] + l[841] + l[847] + l[859] + l[872] + l[878] + l[885] + l[886] + l[888] + l[894] + l[912] + l[915] + l[917] + l[919] + l[925] + l[936] + l[937] + l[950] + l[952] + l[954] + l[956] + l[959] + l[968] + l[970] + l[973] + l[982] + l[984] + l[996] + l[1009] + l[1015] + l[1035] + l[1050] + l[1054] + l[1062] + l[1063] + l[1065] + l[1076] + l[1083] + l[1086] + l[1099] + l[1105] + l[1111] + l[1117] + l[1119] + l[1126] + l[1129] + l[1132] + l[1135] + l[1138] + l[1141] + l[1143] + l[1163] + l[1165] + l[1173] + l[1202] + l[1209] + l[1219] + l[1231] + l[1233] + l[1238] + l[1244] + l[1249] + l[1255] + l[1259] + l[1266] + l[1273] + l[1275] + l[1288] + l[1295] + l[1313] + l[1328] + l[1342] + l[1346] + l[1365] + l[1374]; // 0.125
	assign val[9] = l[7] + l[25] + l[34] + l[36] + l[42] + l[44] + l[47] + l[49] + l[50] + l[52] + l[55] + l[64] + l[77] + l[81] + l[83] + l[88] + l[89] + l[101] + l[112] + l[114] + l[120] + l[122] + l[124] + l[132] + l[135] + l[136] + l[138] + l[141] + l[142] + l[148] + l[165] + l[168] + l[175] + l[176] + l[178] + l[182] + l[187] + l[190] + l[193] + l[197] + l[200] + l[203] + l[206] + l[210] + l[211] + l[216] + l[236] + l[256] + l[259] + l[276] + l[277] + l[286] + l[290] + l[296] + l[309] + l[311] + l[320] + l[326] + l[328] + l[333] + l[339] + l[353] + l[356] + l[364] + l[372] + l[374] + l[379] + l[382] + l[385] + l[401] + l[412] + l[426] + l[429] + l[431] + l[437] + l[460] + l[492] + l[499] + l[520] + l[528] + l[534] + l[545] + l[562] + l[564] + l[593] + l[594] + l[601] + l[603] + l[608] + l[614] + l[635] + l[639] + l[642] + l[645] + l[674] + l[681] + l[691] + l[704] + l[712] + l[713] + l[716] + l[719] + l[721] + l[732] + l[734] + l[765] + l[778] + l[813] + l[829] + l[849] + l[855] + l[892] + l[988] + l[999] + l[1025] + l[1048] + l[1113] + l[1147] + l[1157] + l[1175] + l[1195] + l[1332] + l[1362]; // 0.25
	assign val[10] = l[1] + l[19] + l[20] + l[23] + l[24] + l[30] + l[33] + l[45] + l[58] + l[60] + l[66] + l[70] + l[74] + l[92] + l[105] + l[108] + l[116] + l[127] + l[147] + l[172] + l[231] + l[241] + l[335] + l[373] + l[402] + l[485] + l[519] + l[539] + l[1058]; // 0.5
	assign val[11] = l[4] + l[11] + l[14] + l[69] + l[123] + l[321]; // 1.0
	assign val[12] = l[2] + l[8]; // 2.0
endmodule

module leaf_counter_3(input logic [0:1472] l, output logic [7:0] val [0:12]);
	assign val[0] = l[1] + l[32] + l[70] + l[102] + l[125] + l[149] + l[185] + l[202] + l[218] + l[251] + l[253] + l[263] + l[264] + l[268] + l[282] + l[301] + l[307] + l[311] + l[345] + l[362] + l[364] + l[373] + l[374] + l[386] + l[391] + l[448] + l[477] + l[494] + l[510] + l[541] + l[557] + l[568] + l[612] + l[645] + l[658] + l[661] + l[690] + l[696] + l[741] + l[745] + l[751] + l[790] + l[809] + l[815] + l[829] + l[863] + l[983] + l[987] + l[1000] + l[1014] + l[1060] + l[1102] + l[1120] + l[1153] + l[1200] + l[1253] + l[1263] + l[1280] + l[1410]; // -0.25
	assign val[1] = l[0] + l[2] + l[4] + l[7] + l[13] + l[14] + l[16] + l[19] + l[20] + l[23] + l[26] + l[28] + l[31] + l[33] + l[34] + l[37] + l[38] + l[43] + l[46] + l[51] + l[52] + l[56] + l[57] + l[59] + l[60] + l[63] + l[65] + l[66] + l[68] + l[72] + l[74] + l[76] + l[79] + l[80] + l[85] + l[86] + l[92] + l[95] + l[98] + l[100] + l[103] + l[104] + l[105] + l[107] + l[108] + l[112] + l[114] + l[117] + l[123] + l[127] + l[128] + l[131] + l[136] + l[139] + l[142] + l[146] + l[147] + l[151] + l[155] + l[157] + l[163] + l[166] + l[170] + l[172] + l[175] + l[183] + l[186] + l[188] + l[189] + l[195] + l[199] + l[201] + l[203] + l[206] + l[208] + l[210] + l[212] + l[215] + l[216] + l[221] + l[222] + l[226] + l[228] + l[233] + l[245] + l[247] + l[248] + l[255] + l[260] + l[267] + l[271] + l[272] + l[275] + l[278] + l[281] + l[285] + l[287] + l[299] + l[305] + l[312] + l[314] + l[321] + l[322] + l[325] + l[329] + l[337] + l[338] + l[342] + l[347] + l[349] + l[353] + l[358] + l[383] + l[384] + l[388] + l[389] + l[394] + l[399] + l[401] + l[404] + l[406] + l[407] + l[413] + l[421] + l[427] + l[430] + l[436] + l[437] + l[444] + l[447] + l[450] + l[456] + l[458] + l[461] + l[467] + l[470] + l[476] + l[479] + l[480] + l[483] + l[489] + l[493] + l[498] + l[501] + l[505] + l[508] + l[520] + l[522] + l[525] + l[528] + l[535] + l[552] + l[562] + l[570] + l[576] + l[580] + l[584] + l[592] + l[596] + l[598] + l[601] + l[607] + l[608] + l[615] + l[620] + l[622] + l[623] + l[637] + l[647] + l[650] + l[655] + l[657] + l[659] + l[664] + l[665] + l[668] + l[675] + l[683] + l[686] + l[699] + l[704] + l[708] + l[713] + l[730] + l[731] + l[738] + l[742] + l[749] + l[758] + l[771] + l[774] + l[776] + l[783] + l[786] + l[792] + l[793] + l[798] + l[800] + l[802] + l[804] + l[805] + l[807] + l[810] + l[817] + l[821] + l[828] + l[831] + l[845] + l[848] + l[852] + l[853] + l[857] + l[864] + l[870] + l[872] + l[875] + l[879] + l[883] + l[887] + l[888] + l[893] + l[899] + l[901] + l[905] + l[908] + l[918] + l[922] + l[924] + l[929] + l[932] + l[933] + l[945] + l[953] + l[954] + l[963] + l[966] + l[967] + l[970] + l[971] + l[975] + l[989] + l[991] + l[999] + l[1004] + l[1008] + l[1015] + l[1021] + l[1026] + l[1030] + l[1034] + l[1035] + l[1040] + l[1043] + l[1064] + l[1069] + l[1070] + l[1074] + l[1079] + l[1083] + l[1088] + l[1090] + l[1094] + l[1095] + l[1107] + l[1112] + l[1123] + l[1147] + l[1152] + l[1155] + l[1164] + l[1166] + l[1167] + l[1170] + l[1174] + l[1175] + l[1179] + l[1184] + l[1187] + l[1189] + l[1190] + l[1197] + l[1211] + l[1214] + l[1222] + l[1223] + l[1226] + l[1233] + l[1247] + l[1252] + l[1262] + l[1276] + l[1281] + l[1290] + l[1300] + l[1304] + l[1309] + l[1312] + l[1314] + l[1319] + l[1329] + l[1332] + l[1350] + l[1356] + l[1359] + l[1363] + l[1371] + l[1373] + l[1374] + l[1376] + l[1380] + l[1382] + l[1386] + l[1388] + l[1399] + l[1402] + l[1405] + l[1420] + l[1424] + l[1429] + l[1434] + l[1437] + l[1444] + l[1446] + l[1469]; // -0.125
	assign val[2] = l[11] + l[41] + l[44] + l[55] + l[71] + l[77] + l[83] + l[110] + l[119] + l[137] + l[140] + l[144] + l[150] + l[154] + l[159] + l[162] + l[168] + l[177] + l[191] + l[194] + l[213] + l[225] + l[230] + l[234] + l[238] + l[250] + l[262] + l[283] + l[286] + l[292] + l[295] + l[298] + l[317] + l[318] + l[331] + l[356] + l[368] + l[369] + l[371] + l[376] + l[381] + l[387] + l[398] + l[409] + l[424] + l[439] + l[443] + l[455] + l[495] + l[499] + l[503] + l[507] + l[511] + l[514] + l[526] + l[538] + l[546] + l[549] + l[551] + l[558] + l[561] + l[567] + l[571] + l[573] + l[588] + l[603] + l[611] + l[617] + l[630] + l[633] + l[635] + l[638] + l[640] + l[641] + l[648] + l[662] + l[670] + l[682] + l[685] + l[711] + l[716] + l[718] + l[720] + l[725] + l[736] + l[754] + l[764] + l[768] + l[781] + l[811] + l[837] + l[839] + l[860] + l[910] + l[912] + l[920] + l[930] + l[936] + l[942] + l[943] + l[946] + l[947] + l[958] + l[978] + l[979] + l[986] + l[993] + l[995] + l[1010] + l[1018] + l[1031] + l[1042] + l[1045] + l[1050] + l[1051] + l[1054] + l[1061] + l[1062] + l[1089] + l[1092] + l[1105] + l[1106] + l[1115] + l[1126] + l[1136] + l[1162] + l[1178] + l[1193] + l[1194] + l[1207] + l[1213] + l[1215] + l[1217] + l[1219] + l[1229] + l[1230] + l[1234] + l[1239] + l[1245] + l[1249] + l[1250] + l[1256] + l[1257] + l[1264] + l[1265] + l[1283] + l[1285] + l[1289] + l[1292] + l[1298] + l[1305] + l[1316] + l[1325] + l[1334] + l[1337] + l[1338] + l[1340] + l[1343] + l[1347] + l[1355] + l[1360] + l[1365] + l[1394] + l[1397] + l[1412] + l[1426] + l[1442] + l[1451] + l[1453] + l[1456] + l[1457] + l[1460] + l[1465] + l[1472]; // -0.0625
	assign val[3] = l[47] + l[53] + l[88] + l[120] + l[179] + l[217] + l[288] + l[290] + l[302] + l[357] + l[363] + l[365] + l[378] + l[396] + l[405] + l[429] + l[453] + l[462] + l[466] + l[484] + l[542] + l[556] + l[600] + l[627] + l[632] + l[688] + l[692] + l[697] + l[728] + l[744] + l[747] + l[752] + l[765] + l[777] + l[825] + l[841] + l[844] + l[854] + l[862] + l[881] + l[890] + l[892] + l[894] + l[896] + l[915] + l[917] + l[923] + l[938] + l[956] + l[961] + l[1005] + l[1033] + l[1036] + l[1058] + l[1066] + l[1081] + l[1100] + l[1108] + l[1111] + l[1119] + l[1121] + l[1129] + l[1130] + l[1133] + l[1141] + l[1154] + l[1181] + l[1183] + l[1202] + l[1221] + l[1232] + l[1236] + l[1240] + l[1242] + l[1254] + l[1272] + l[1287] + l[1291] + l[1311] + l[1326] + l[1358] + l[1362] + l[1364] + l[1378] + l[1381] + l[1389] + l[1403] + l[1406] + l[1414] + l[1423] + l[1436] + l[1440] + l[1447] + l[1463]; // -0.03125
	assign val[4] = l[124] + l[197] + l[200] + l[254] + l[326] + l[334] + l[411] + l[529] + l[544] + l[565] + l[578] + l[606] + l[680] + l[719] + l[724] + l[733] + l[772] + l[787] + l[789] + l[806] + l[867] + l[884] + l[964] + l[976] + l[997] + l[1006] + l[1016] + l[1019] + l[1024] + l[1038] + l[1057] + l[1065] + l[1077] + l[1078] + l[1097] + l[1103] + l[1140] + l[1160] + l[1168] + l[1185] + l[1205] + l[1259] + l[1277] + l[1279] + l[1299] + l[1303] + l[1313] + l[1318] + l[1321] + l[1353] + l[1367] + l[1396] + l[1431] + l[1449]; // -0.015625
	assign val[5] = l[97] + l[176] + l[229] + l[360] + l[425] + l[438] + l[457] + l[515] + l[553] + l[569] + l[581] + l[643] + l[654] + l[663] + l[666] + l[693] + l[710] + l[735] + l[753] + l[759] + l[763] + l[775] + l[794] + l[795] + l[797] + l[885] + l[906] + l[941] + l[944] + l[977] + l[1027] + l[1046] + l[1068] + l[1104] + l[1109] + l[1145] + l[1151] + l[1173] + l[1180] + l[1196] + l[1203] + l[1210] + l[1243] + l[1275] + l[1295] + l[1315] + l[1352] + l[1379] + l[1385] + l[1445] + l[1462]; // 0.015625
	assign val[6] = l[25] + l[50] + l[129] + l[152] + l[182] + l[190] + l[237] + l[239] + l[243] + l[244] + l[257] + l[273] + l[279] + l[297] + l[336] + l[350] + l[351] + l[419] + l[422] + l[428] + l[451] + l[454] + l[524] + l[534] + l[560] + l[597] + l[624] + l[625] + l[660] + l[694] + l[732] + l[739] + l[762] + l[816] + l[847] + l[858] + l[880] + l[898] + l[900] + l[919] + l[952] + l[960] + l[968] + l[980] + l[994] + l[1022] + l[1025] + l[1029] + l[1044] + l[1052] + l[1067] + l[1071] + l[1156] + l[1169] + l[1171] + l[1199] + l[1209] + l[1227] + l[1235] + l[1261] + l[1297] + l[1310] + l[1327] + l[1328] + l[1330] + l[1333] + l[1335] + l[1341] + l[1369] + l[1383] + l[1391] + l[1398] + l[1401] + l[1409] + l[1415] + l[1416] + l[1425] + l[1427] + l[1432] + l[1435] + l[1452]; // 0.03125
	assign val[7] = l[21] + l[106] + l[130] + l[156] + l[158] + l[171] + l[209] + l[211] + l[227] + l[240] + l[246] + l[249] + l[261] + l[269] + l[270] + l[284] + l[294] + l[300] + l[303] + l[306] + l[309] + l[310] + l[320] + l[335] + l[339] + l[343] + l[344] + l[355] + l[361] + l[366] + l[375] + l[379] + l[390] + l[395] + l[400] + l[403] + l[412] + l[414] + l[441] + l[445] + l[446] + l[449] + l[472] + l[485] + l[487] + l[491] + l[500] + l[502] + l[506] + l[509] + l[518] + l[547] + l[548] + l[564] + l[575] + l[577] + l[586] + l[589] + l[595] + l[599] + l[602] + l[605] + l[614] + l[619] + l[629] + l[634] + l[642] + l[644] + l[649] + l[653] + l[667] + l[681] + l[684] + l[687] + l[707] + l[712] + l[714] + l[715] + l[723] + l[726] + l[734] + l[767] + l[780] + l[784] + l[799] + l[803] + l[822] + l[824] + l[827] + l[846] + l[856] + l[871] + l[873] + l[874] + l[882] + l[886] + l[889] + l[897] + l[902] + l[909] + l[911] + l[914] + l[921] + l[925] + l[926] + l[937] + l[957] + l[962] + l[988] + l[1007] + l[1011] + l[1023] + l[1041] + l[1047] + l[1049] + l[1053] + l[1055] + l[1059] + l[1073] + l[1075] + l[1085] + l[1093] + l[1113] + l[1117] + l[1122] + l[1134] + l[1137] + l[1138] + l[1163] + l[1165] + l[1177] + l[1192] + l[1204] + l[1206] + l[1212] + l[1224] + l[1238] + l[1244] + l[1246] + l[1270] + l[1271] + l[1274] + l[1282] + l[1286] + l[1288] + l[1293] + l[1296] + l[1322] + l[1339] + l[1372] + l[1393] + l[1395] + l[1404] + l[1439] + l[1450] + l[1454] + l[1459] + l[1466] + l[1471]; // 0.0625
	assign val[8] = l[39] + l[42] + l[69] + l[84] + l[89] + l[99] + l[111] + l[135] + l[141] + l[143] + l[145] + l[148] + l[153] + l[160] + l[161] + l[167] + l[169] + l[180] + l[184] + l[192] + l[193] + l[204] + l[207] + l[220] + l[223] + l[224] + l[231] + l[232] + l[235] + l[236] + l[242] + l[252] + l[259] + l[266] + l[274] + l[276] + l[291] + l[293] + l[296] + l[304] + l[315] + l[316] + l[323] + l[327] + l[328] + l[340] + l[348] + l[352] + l[367] + l[370] + l[377] + l[380] + l[382] + l[415] + l[417] + l[426] + l[435] + l[459] + l[460] + l[469] + l[478] + l[482] + l[488] + l[512] + l[519] + l[521] + l[530] + l[537] + l[540] + l[543] + l[545] + l[550] + l[559] + l[591] + l[593] + l[618] + l[626] + l[628] + l[631] + l[639] + l[646] + l[651] + l[656] + l[672] + l[673] + l[676] + l[678] + l[679] + l[691] + l[698] + l[702] + l[706] + l[717] + l[721] + l[729] + l[746] + l[755] + l[760] + l[766] + l[769] + l[773] + l[778] + l[788] + l[796] + l[808] + l[814] + l[818] + l[826] + l[832] + l[835] + l[838] + l[851] + l[861] + l[866] + l[869] + l[876] + l[891] + l[895] + l[907] + l[913] + l[916] + l[931] + l[935] + l[948] + l[951] + l[965] + l[969] + l[974] + l[996] + l[1003] + l[1017] + l[1020] + l[1028] + l[1032] + l[1048] + l[1063] + l[1080] + l[1084] + l[1087] + l[1091] + l[1099] + l[1101] + l[1118] + l[1124] + l[1127] + l[1128] + l[1131] + l[1144] + l[1146] + l[1150] + l[1158] + l[1159] + l[1161] + l[1172] + l[1182] + l[1186] + l[1198] + l[1201] + l[1216] + l[1220] + l[1225] + l[1228] + l[1231] + l[1237] + l[1241] + l[1248] + l[1251] + l[1255] + l[1260] + l[1268] + l[1278] + l[1302] + l[1306] + l[1307] + l[1317] + l[1320] + l[1324] + l[1331] + l[1336] + l[1344] + l[1346] + l[1348] + l[1351] + l[1354] + l[1357] + l[1368] + l[1377] + l[1390] + l[1392] + l[1400] + l[1407] + l[1413] + l[1417] + l[1418] + l[1428] + l[1448] + l[1455] + l[1461] + l[1464] + l[1467]; // 0.125
	assign val[9] = l[15] + l[17] + l[18] + l[27] + l[29] + l[35] + l[36] + l[45] + l[48] + l[58] + l[61] + l[62] + l[64] + l[67] + l[75] + l[78] + l[81] + l[90] + l[93] + l[94] + l[96] + l[101] + l[109] + l[113] + l[115] + l[118] + l[121] + l[122] + l[126] + l[138] + l[164] + l[165] + l[173] + l[178] + l[181] + l[187] + l[198] + l[205] + l[214] + l[241] + l[256] + l[277] + l[280] + l[289] + l[308] + l[313] + l[319] + l[324] + l[330] + l[341] + l[354] + l[359] + l[385] + l[397] + l[416] + l[420] + l[423] + l[432] + l[434] + l[442] + l[452] + l[463] + l[464] + l[471] + l[474] + l[490] + l[497] + l[516] + l[517] + l[527] + l[532] + l[533] + l[555] + l[566] + l[572] + l[574] + l[582] + l[587] + l[616] + l[636] + l[669] + l[689] + l[695] + l[701] + l[709] + l[727] + l[740] + l[750] + l[756] + l[761] + l[782] + l[785] + l[801] + l[833] + l[842] + l[843] + l[849] + l[878] + l[903] + l[927] + l[939] + l[949] + l[959] + l[981] + l[985] + l[992] + l[1012] + l[1037] + l[1056] + l[1076] + l[1086] + l[1110] + l[1114] + l[1125] + l[1132] + l[1139] + l[1195] + l[1208] + l[1294] + l[1361] + l[1370] + l[1384]; // 0.25
	assign val[10] = l[3] + l[5] + l[6] + l[8] + l[10] + l[12] + l[22] + l[24] + l[30] + l[40] + l[54] + l[82] + l[87] + l[132] + l[219] + l[333] + l[372] + l[408] + l[418] + l[433] + l[523] + l[539] + l[585] + l[594] + l[610] + l[674] + l[819] + l[836] + l[1072]; // 0.5
	assign val[11] = l[9] + l[134] + l[332]; // 1.0
	assign val[12] = 0; // 2.0
endmodule

module leaf_counter_4(input logic [0:1315] l, output logic [7:0] val [0:12]);
	assign val[0] = l[8] + l[11] + l[16] + l[27] + l[29] + l[36] + l[47] + l[60] + l[69] + l[73] + l[79] + l[81] + l[86] + l[91] + l[103] + l[106] + l[140] + l[148] + l[162] + l[164] + l[170] + l[180] + l[216] + l[226] + l[234] + l[265] + l[270] + l[272] + l[280] + l[290] + l[296] + l[300] + l[309] + l[316] + l[327] + l[329] + l[332] + l[337] + l[345] + l[367] + l[383] + l[392] + l[413] + l[420] + l[422] + l[423] + l[426] + l[443] + l[447] + l[449] + l[450] + l[462] + l[485] + l[486] + l[494] + l[519] + l[529] + l[531] + l[532] + l[535] + l[538] + l[547] + l[549] + l[556] + l[557] + l[568] + l[580] + l[591] + l[593] + l[603] + l[621] + l[622] + l[631] + l[632] + l[640] + l[643] + l[645] + l[670] + l[687] + l[695] + l[698] + l[704] + l[717] + l[731] + l[740] + l[744] + l[759] + l[782] + l[794] + l[816] + l[822] + l[834] + l[846] + l[862] + l[892] + l[899] + l[902] + l[906] + l[919] + l[926] + l[940] + l[956] + l[986] + l[993] + l[1007] + l[1048] + l[1058] + l[1254]; // -0.25
	assign val[1] = l[0] + l[3] + l[6] + l[9] + l[10] + l[13] + l[15] + l[17] + l[18] + l[21] + l[23] + l[28] + l[32] + l[35] + l[37] + l[39] + l[40] + l[45] + l[46] + l[48] + l[51] + l[52] + l[57] + l[63] + l[66] + l[68] + l[72] + l[75] + l[77] + l[80] + l[83] + l[84] + l[94] + l[96] + l[99] + l[104] + l[109] + l[111] + l[113] + l[114] + l[116] + l[117] + l[119] + l[121] + l[123] + l[124] + l[127] + l[129] + l[131] + l[136] + l[139] + l[142] + l[145] + l[146] + l[149] + l[151] + l[153] + l[154] + l[156] + l[159] + l[161] + l[163] + l[165] + l[167] + l[172] + l[175] + l[177] + l[178] + l[181] + l[183] + l[184] + l[187] + l[191] + l[192] + l[195] + l[196] + l[198] + l[203] + l[207] + l[208] + l[211] + l[214] + l[218] + l[221] + l[222] + l[223] + l[230] + l[232] + l[235] + l[238] + l[239] + l[241] + l[246] + l[247] + l[252] + l[253] + l[256] + l[259] + l[261] + l[264] + l[267] + l[269] + l[274] + l[284] + l[287] + l[289] + l[292] + l[295] + l[298] + l[303] + l[304] + l[310] + l[312] + l[314] + l[319] + l[320] + l[324] + l[330] + l[336] + l[344] + l[346] + l[348] + l[350] + l[353] + l[356] + l[358] + l[360] + l[361] + l[364] + l[371] + l[373] + l[376] + l[381] + l[386] + l[388] + l[393] + l[396] + l[398] + l[400] + l[404] + l[406] + l[416] + l[418] + l[425] + l[427] + l[430] + l[432] + l[433] + l[437] + l[451] + l[452] + l[454] + l[465] + l[469] + l[470] + l[475] + l[476] + l[478] + l[481] + l[483] + l[487] + l[489] + l[490] + l[492] + l[495] + l[498] + l[501] + l[503] + l[512] + l[514] + l[521] + l[524] + l[537] + l[539] + l[544] + l[546] + l[554] + l[562] + l[570] + l[572] + l[573] + l[576] + l[578] + l[587] + l[597] + l[600] + l[605] + l[608] + l[613] + l[615] + l[616] + l[625] + l[629] + l[635] + l[637] + l[642] + l[648] + l[651] + l[656] + l[660] + l[665] + l[667] + l[675] + l[678] + l[681] + l[686] + l[688] + l[692] + l[700] + l[702] + l[705] + l[714] + l[715] + l[721] + l[726] + l[739] + l[743] + l[745] + l[747] + l[748] + l[751] + l[752] + l[753] + l[756] + l[765] + l[768] + l[773] + l[779] + l[781] + l[787] + l[788] + l[791] + l[798] + l[804] + l[809] + l[811] + l[817] + l[830] + l[833] + l[839] + l[843] + l[845] + l[850] + l[854] + l[856] + l[859] + l[861] + l[869] + l[873] + l[874] + l[878] + l[881] + l[882] + l[896] + l[897] + l[904] + l[910] + l[911] + l[913] + l[915] + l[917] + l[920] + l[925] + l[929] + l[931] + l[936] + l[939] + l[942] + l[948] + l[949] + l[950] + l[955] + l[959] + l[964] + l[969] + l[972] + l[973] + l[978] + l[985] + l[987] + l[990] + l[991] + l[1001] + l[1009] + l[1011] + l[1013] + l[1015] + l[1023] + l[1024] + l[1025] + l[1028] + l[1031] + l[1034] + l[1038] + l[1040] + l[1042] + l[1046] + l[1056] + l[1071] + l[1073] + l[1074] + l[1077] + l[1083] + l[1086] + l[1091] + l[1096] + l[1101] + l[1104] + l[1105] + l[1106] + l[1108] + l[1114] + l[1121] + l[1127] + l[1129] + l[1133] + l[1138] + l[1140] + l[1141] + l[1148] + l[1152] + l[1155] + l[1157] + l[1160] + l[1161] + l[1172] + l[1173] + l[1176] + l[1185] + l[1189] + l[1196] + l[1197] + l[1201] + l[1203] + l[1206] + l[1208] + l[1212] + l[1215] + l[1216] + l[1219] + l[1230] + l[1237] + l[1238] + l[1243] + l[1244] + l[1247] + l[1255] + l[1261] + l[1266] + l[1267] + l[1270] + l[1272] + l[1276] + l[1279] + l[1281] + l[1287] + l[1294] + l[1306] + l[1314] + l[1315]; // -0.125
	assign val[2] = l[31] + l[43] + l[55] + l[65] + l[87] + l[92] + l[101] + l[107] + l[125] + l[133] + l[137] + l[141] + l[147] + l[171] + l[179] + l[205] + l[213] + l[217] + l[219] + l[228] + l[262] + l[271] + l[273] + l[278] + l[283] + l[293] + l[301] + l[328] + l[334] + l[340] + l[341] + l[362] + l[370] + l[378] + l[380] + l[390] + l[391] + l[405] + l[409] + l[414] + l[419] + l[421] + l[428] + l[435] + l[439] + l[444] + l[448] + l[461] + l[463] + l[497] + l[509] + l[511] + l[523] + l[527] + l[528] + l[533] + l[534] + l[540] + l[548] + l[555] + l[558] + l[561] + l[564] + l[574] + l[582] + l[592] + l[594] + l[595] + l[602] + l[607] + l[623] + l[633] + l[661] + l[664] + l[671] + l[677] + l[682] + l[690] + l[693] + l[696] + l[707] + l[710] + l[719] + l[729] + l[736] + l[741] + l[750] + l[760] + l[764] + l[771] + l[793] + l[795] + l[800] + l[814] + l[821] + l[823] + l[826] + l[829] + l[837] + l[847] + l[853] + l[863] + l[871] + l[891] + l[893] + l[898] + l[907] + l[912] + l[951] + l[996] + l[1005] + l[1008] + l[1016] + l[1035] + l[1041] + l[1050] + l[1053] + l[1060] + l[1064] + l[1067] + l[1078] + l[1117] + l[1120] + l[1135] + l[1150] + l[1164] + l[1167] + l[1170] + l[1178] + l[1183] + l[1187] + l[1192] + l[1217] + l[1222] + l[1226] + l[1232] + l[1245] + l[1253] + l[1262] + l[1291] + l[1295] + l[1298]; // -0.0625
	assign val[3] = l[22] + l[70] + l[105] + l[115] + l[157] + l[201] + l[202] + l[225] + l[236] + l[281] + l[297] + l[366] + l[399] + l[411] + l[441] + l[455] + l[457] + l[459] + l[466] + l[515] + l[542] + l[559] + l[579] + l[584] + l[585] + l[610] + l[620] + l[626] + l[649] + l[655] + l[697] + l[718] + l[722] + l[724] + l[732] + l[734] + l[785] + l[803] + l[819] + l[824] + l[835] + l[844] + l[865] + l[866] + l[868] + l[886] + l[894] + l[945] + l[953] + l[957] + l[968] + l[975] + l[982] + l[1027] + l[1033] + l[1055] + l[1059] + l[1063] + l[1069] + l[1072] + l[1093] + l[1100] + l[1107] + l[1110] + l[1125] + l[1146] + l[1168] + l[1194] + l[1200] + l[1202] + l[1207] + l[1209] + l[1235] + l[1251] + l[1268] + l[1283] + l[1307] + l[1312]; // -0.03125
	assign val[4] = l[41] + l[78] + l[89] + l[97] + l[242] + l[244] + l[254] + l[277] + l[291] + l[315] + l[317] + l[384] + l[464] + l[506] + l[612] + l[630] + l[639] + l[666] + l[669] + l[679] + l[706] + l[712] + l[813] + l[842] + l[849] + l[888] + l[901] + l[916] + l[927] + l[946] + l[962] + l[963] + l[966] + l[1018] + l[1021] + l[1029] + l[1047] + l[1111] + l[1180] + l[1225] + l[1228] + l[1240] + l[1264] + l[1274] + l[1282] + l[1285] + l[1301]; // -0.015625
	assign val[5] = l[49] + l[85] + l[130] + l[190] + l[199] + l[311] + l[321] + l[326] + l[349] + l[352] + l[375] + l[440] + l[474] + l[518] + l[525] + l[604] + l[627] + l[636] + l[647] + l[650] + l[709] + l[725] + l[783] + l[792] + l[801] + l[851] + l[872] + l[876] + l[880] + l[883] + l[884] + l[900] + l[924] + l[932] + l[943] + l[947] + l[954] + l[960] + l[970] + l[992] + l[1019] + l[1043] + l[1061] + l[1103] + l[1109] + l[1122] + l[1147] + l[1156] + l[1162] + l[1169] + l[1179] + l[1186] + l[1277] + l[1288] + l[1309]; // 0.015625
	assign val[6] = l[50] + l[53] + l[61] + l[110] + l[120] + l[168] + l[185] + l[189] + l[249] + l[266] + l[307] + l[308] + l[347] + l[395] + l[397] + l[401] + l[415] + l[429] + l[480] + l[484] + l[499] + l[516] + l[520] + l[543] + l[553] + l[571] + l[577] + l[581] + l[601] + l[609] + l[614] + l[617] + l[619] + l[628] + l[663] + l[672] + l[674] + l[685] + l[735] + l[742] + l[754] + l[758] + l[766] + l[799] + l[802] + l[818] + l[827] + l[836] + l[858] + l[860] + l[875] + l[890] + l[909] + l[914] + l[921] + l[928] + l[952] + l[967] + l[980] + l[984] + l[997] + l[1012] + l[1026] + l[1030] + l[1045] + l[1052] + l[1054] + l[1092] + l[1097] + l[1139] + l[1184] + l[1188] + l[1190] + l[1199] + l[1210] + l[1223] + l[1246] + l[1265] + l[1269] + l[1280] + l[1293] + l[1296] + l[1305] + l[1311]; // 0.03125
	assign val[7] = l[1] + l[25] + l[56] + l[62] + l[90] + l[112] + l[134] + l[144] + l[155] + l[160] + l[176] + l[186] + l[194] + l[206] + l[210] + l[215] + l[224] + l[245] + l[248] + l[255] + l[257] + l[260] + l[268] + l[276] + l[286] + l[294] + l[299] + l[302] + l[313] + l[318] + l[357] + l[363] + l[369] + l[377] + l[387] + l[389] + l[394] + l[403] + l[410] + l[412] + l[431] + l[442] + l[445] + l[456] + l[458] + l[460] + l[468] + l[471] + l[493] + l[496] + l[505] + l[510] + l[541] + l[560] + l[565] + l[569] + l[583] + l[586] + l[588] + l[590] + l[596] + l[599] + l[611] + l[634] + l[644] + l[662] + l[680] + l[683] + l[691] + l[708] + l[711] + l[716] + l[727] + l[733] + l[737] + l[738] + l[749] + l[755] + l[763] + l[767] + l[775] + l[780] + l[789] + l[805] + l[807] + l[820] + l[832] + l[848] + l[857] + l[867] + l[879] + l[918] + l[937] + l[938] + l[958] + l[979] + l[995] + l[1003] + l[1014] + l[1020] + l[1022] + l[1032] + l[1036] + l[1039] + l[1049] + l[1057] + l[1062] + l[1065] + l[1075] + l[1076] + l[1079] + l[1087] + l[1112] + l[1115] + l[1118] + l[1119] + l[1124] + l[1126] + l[1142] + l[1143] + l[1149] + l[1153] + l[1159] + l[1163] + l[1165] + l[1166] + l[1181] + l[1182] + l[1195] + l[1213] + l[1221] + l[1229] + l[1231] + l[1233] + l[1234] + l[1239] + l[1249] + l[1252] + l[1257] + l[1273] + l[1284] + l[1300] + l[1304] + l[1308]; // 0.0625
	assign val[8] = l[5] + l[33] + l[38] + l[44] + l[59] + l[82] + l[95] + l[98] + l[100] + l[122] + l[128] + l[132] + l[150] + l[152] + l[166] + l[169] + l[173] + l[182] + l[188] + l[193] + l[197] + l[200] + l[204] + l[212] + l[220] + l[227] + l[229] + l[233] + l[243] + l[251] + l[258] + l[279] + l[282] + l[288] + l[306] + l[322] + l[325] + l[333] + l[335] + l[339] + l[343] + l[351] + l[355] + l[365] + l[372] + l[379] + l[382] + l[385] + l[402] + l[436] + l[438] + l[446] + l[453] + l[467] + l[473] + l[477] + l[479] + l[500] + l[507] + l[517] + l[526] + l[536] + l[545] + l[552] + l[575] + l[598] + l[606] + l[618] + l[624] + l[641] + l[657] + l[659] + l[689] + l[694] + l[699] + l[720] + l[723] + l[761] + l[770] + l[772] + l[777] + l[778] + l[784] + l[790] + l[797] + l[806] + l[812] + l[825] + l[828] + l[831] + l[838] + l[855] + l[864] + l[885] + l[887] + l[889] + l[895] + l[923] + l[934] + l[961] + l[965] + l[983] + l[999] + l[1002] + l[1006] + l[1017] + l[1037] + l[1044] + l[1051] + l[1066] + l[1068] + l[1070] + l[1081] + l[1085] + l[1088] + l[1094] + l[1099] + l[1145] + l[1154] + l[1171] + l[1177] + l[1193] + l[1224] + l[1227] + l[1236] + l[1241] + l[1250] + l[1278] + l[1286] + l[1289] + l[1292] + l[1297] + l[1310]; // 0.125
	assign val[9] = l[20] + l[54] + l[58] + l[64] + l[67] + l[71] + l[74] + l[76] + l[88] + l[93] + l[102] + l[108] + l[118] + l[126] + l[135] + l[138] + l[158] + l[174] + l[250] + l[263] + l[408] + l[488] + l[522] + l[638] + l[653] + l[658] + l[668] + l[701] + l[713] + l[730] + l[757] + l[808] + l[841] + l[852] + l[870] + l[877] + l[935] + l[944] + l[977] + l[981] + l[998] + l[1082] + l[1116] + l[1131] + l[1137] + l[1144] + l[1191] + l[1205] + l[1259] + l[1303]; // 0.25
	assign val[10] = l[2] + l[12] + l[19] + l[24] + l[30] + l[34] + l[42] + l[933]; // 0.5
	assign val[11] = l[4] + l[7]; // 1.0
	assign val[12] = 0; // 2.0
endmodule

module leaf_counter_5(input logic [0:1401] l, output logic [7:0] val [0:12]);
	assign val[0] = l[5] + l[7] + l[10] + l[14] + l[20] + l[21] + l[32] + l[37] + l[38] + l[44] + l[49] + l[56] + l[59] + l[60] + l[85] + l[87] + l[104] + l[106] + l[124] + l[131] + l[149] + l[152] + l[154] + l[172] + l[179] + l[180] + l[184] + l[186] + l[192] + l[240] + l[242] + l[263] + l[273] + l[278] + l[312] + l[315] + l[348] + l[362] + l[370] + l[379] + l[386] + l[442] + l[461] + l[517] + l[528] + l[529] + l[537] + l[540] + l[541] + l[544] + l[553] + l[594] + l[601] + l[603] + l[607] + l[628] + l[650] + l[681] + l[700] + l[715] + l[726] + l[732] + l[742] + l[770] + l[792] + l[798] + l[802] + l[803] + l[836] + l[837] + l[839] + l[852] + l[863] + l[867] + l[883] + l[962] + l[969] + l[987] + l[1014] + l[1023] + l[1060] + l[1121] + l[1201] + l[1212] + l[1238] + l[1262] + l[1281] + l[1331]; // -0.25
	assign val[1] = l[0] + l[13] + l[15] + l[18] + l[23] + l[24] + l[28] + l[34] + l[41] + l[48] + l[50] + l[53] + l[55] + l[62] + l[65] + l[69] + l[71] + l[72] + l[75] + l[77] + l[79] + l[80] + l[82] + l[86] + l[89] + l[92] + l[95] + l[96] + l[98] + l[101] + l[103] + l[105] + l[109] + l[112] + l[113] + l[114] + l[119] + l[121] + l[122] + l[129] + l[132] + l[136] + l[138] + l[140] + l[141] + l[143] + l[144] + l[146] + l[153] + l[155] + l[157] + l[160] + l[165] + l[166] + l[169] + l[176] + l[188] + l[194] + l[195] + l[200] + l[202] + l[203] + l[210] + l[212] + l[214] + l[216] + l[219] + l[224] + l[226] + l[228] + l[233] + l[235] + l[236] + l[243] + l[247] + l[249] + l[252] + l[256] + l[259] + l[264] + l[265] + l[271] + l[274] + l[280] + l[282] + l[287] + l[289] + l[291] + l[294] + l[296] + l[300] + l[308] + l[311] + l[314] + l[320] + l[325] + l[332] + l[337] + l[339] + l[340] + l[342] + l[344] + l[347] + l[355] + l[356] + l[358] + l[365] + l[366] + l[371] + l[372] + l[374] + l[382] + l[388] + l[389] + l[395] + l[398] + l[409] + l[412] + l[416] + l[419] + l[420] + l[425] + l[427] + l[432] + l[440] + l[444] + l[448] + l[450] + l[451] + l[456] + l[458] + l[464] + l[465] + l[473] + l[475] + l[481] + l[486] + l[499] + l[500] + l[502] + l[506] + l[509] + l[515] + l[526] + l[533] + l[536] + l[545] + l[560] + l[567] + l[569] + l[575] + l[578] + l[584] + l[587] + l[590] + l[592] + l[599] + l[615] + l[620] + l[633] + l[635] + l[637] + l[639] + l[649] + l[652] + l[655] + l[662] + l[677] + l[679] + l[682] + l[684] + l[690] + l[698] + l[702] + l[705] + l[706] + l[708] + l[712] + l[718] + l[723] + l[728] + l[739] + l[746] + l[753] + l[755] + l[758] + l[761] + l[762] + l[765] + l[769] + l[778] + l[779] + l[784] + l[787] + l[790] + l[795] + l[811] + l[815] + l[816] + l[819] + l[821] + l[831] + l[832] + l[842] + l[848] + l[855] + l[864] + l[879] + l[892] + l[893] + l[898] + l[900] + l[906] + l[913] + l[914] + l[917] + l[919] + l[942] + l[947] + l[951] + l[953] + l[966] + l[975] + l[976] + l[978] + l[985] + l[988] + l[996] + l[1002] + l[1013] + l[1022] + l[1025] + l[1036] + l[1048] + l[1052] + l[1055] + l[1067] + l[1075] + l[1080] + l[1083] + l[1087] + l[1092] + l[1093] + l[1101] + l[1106] + l[1109] + l[1116] + l[1127] + l[1130] + l[1133] + l[1135] + l[1145] + l[1147] + l[1153] + l[1161] + l[1165] + l[1168] + l[1176] + l[1178] + l[1186] + l[1187] + l[1196] + l[1197] + l[1203] + l[1223] + l[1228] + l[1230] + l[1235] + l[1244] + l[1245] + l[1254] + l[1258] + l[1268] + l[1269] + l[1278] + l[1292] + l[1295] + l[1303] + l[1305] + l[1313] + l[1321] + l[1328] + l[1337] + l[1339] + l[1345] + l[1348] + l[1354] + l[1356] + l[1370] + l[1371] + l[1377] + l[1378] + l[1386] + l[1394] + l[1395] + l[1401]; // -0.125
	assign val[2] = l[11] + l[27] + l[45] + l[61] + l[126] + l[134] + l[151] + l[159] + l[173] + l[175] + l[183] + l[185] + l[190] + l[205] + l[209] + l[229] + l[232] + l[237] + l[248] + l[250] + l[262] + l[279] + l[290] + l[297] + l[301] + l[304] + l[317] + l[378] + l[387] + l[391] + l[400] + l[407] + l[436] + l[452] + l[453] + l[470] + l[487] + l[497] + l[519] + l[559] + l[564] + l[565] + l[580] + l[593] + l[597] + l[602] + l[606] + l[612] + l[617] + l[641] + l[645] + l[656] + l[659] + l[665] + l[668] + l[673] + l[675] + l[693] + l[695] + l[710] + l[725] + l[733] + l[734] + l[737] + l[757] + l[767] + l[775] + l[782] + l[800] + l[806] + l[824] + l[827] + l[828] + l[857] + l[859] + l[861] + l[868] + l[871] + l[877] + l[889] + l[890] + l[894] + l[903] + l[909] + l[927] + l[931] + l[937] + l[941] + l[954] + l[957] + l[961] + l[973] + l[993] + l[1000] + l[1003] + l[1006] + l[1015] + l[1020] + l[1024] + l[1027] + l[1039] + l[1041] + l[1046] + l[1049] + l[1050] + l[1064] + l[1069] + l[1098] + l[1118] + l[1136] + l[1138] + l[1143] + l[1154] + l[1155] + l[1157] + l[1160] + l[1170] + l[1208] + l[1218] + l[1221] + l[1226] + l[1237] + l[1247] + l[1249] + l[1272] + l[1274] + l[1275] + l[1284] + l[1286] + l[1288] + l[1298] + l[1300] + l[1307] + l[1311] + l[1316] + l[1322] + l[1330] + l[1332] + l[1336] + l[1340] + l[1341] + l[1344] + l[1359] + l[1361] + l[1375] + l[1385] + l[1389] + l[1392] + l[1399]; // -0.0625
	assign val[3] = l[16] + l[67] + l[117] + l[204] + l[207] + l[218] + l[254] + l[257] + l[266] + l[275] + l[281] + l[299] + l[309] + l[313] + l[327] + l[373] + l[392] + l[411] + l[414] + l[429] + l[446] + l[462] + l[466] + l[468] + l[471] + l[490] + l[492] + l[511] + l[514] + l[522] + l[530] + l[531] + l[534] + l[547] + l[549] + l[568] + l[586] + l[613] + l[616] + l[621] + l[638] + l[647] + l[660] + l[666] + l[687] + l[697] + l[701] + l[709] + l[717] + l[736] + l[747] + l[749] + l[752] + l[763] + l[777] + l[807] + l[810] + l[822] + l[840] + l[845] + l[849] + l[850] + l[866] + l[874] + l[876] + l[887] + l[904] + l[916] + l[936] + l[945] + l[948] + l[952] + l[958] + l[979] + l[982] + l[994] + l[998] + l[1004] + l[1009] + l[1010] + l[1018] + l[1029] + l[1053] + l[1061] + l[1072] + l[1074] + l[1082] + l[1090] + l[1094] + l[1096] + l[1103] + l[1105] + l[1113] + l[1124] + l[1129] + l[1132] + l[1150] + l[1162] + l[1163] + l[1172] + l[1180] + l[1191] + l[1199] + l[1207] + l[1216] + l[1232] + l[1264] + l[1266] + l[1270] + l[1279] + l[1289] + l[1318] + l[1358] + l[1368] + l[1379] + l[1380] + l[1382]; // -0.03125
	assign val[4] = l[91] + l[125] + l[215] + l[221] + l[246] + l[284] + l[321] + l[324] + l[351] + l[368] + l[376] + l[384] + l[402] + l[501] + l[561] + l[576] + l[579] + l[623] + l[625] + l[627] + l[631] + l[654] + l[663] + l[688] + l[729] + l[812] + l[846] + l[896] + l[925] + l[933] + l[983] + l[991] + l[1033] + l[1085] + l[1111] + l[1152] + l[1183] + l[1194] + l[1205] + l[1213] + l[1260] + l[1277] + l[1291] + l[1309] + l[1349] + l[1396]; // -0.015625
	assign val[5] = l[1] + l[329] + l[331] + l[336] + l[352] + l[408] + l[431] + l[447] + l[489] + l[498] + l[510] + l[551] + l[554] + l[572] + l[644] + l[653] + l[713] + l[760] + l[785] + l[799] + l[833] + l[872] + l[974] + l[1021] + l[1028] + l[1032] + l[1037] + l[1047] + l[1091] + l[1125] + l[1146] + l[1222] + l[1252] + l[1317] + l[1326] + l[1335] + l[1365] + l[1384] + l[1400]; // 0.015625
	assign val[6] = l[3] + l[57] + l[68] + l[76] + l[93] + l[110] + l[118] + l[189] + l[201] + l[227] + l[268] + l[270] + l[288] + l[307] + l[354] + l[360] + l[405] + l[421] + l[424] + l[433] + l[439] + l[449] + l[463] + l[491] + l[505] + l[585] + l[588] + l[589] + l[611] + l[630] + l[640] + l[669] + l[672] + l[680] + l[691] + l[699] + l[727] + l[735] + l[738] + l[748] + l[750] + l[780] + l[791] + l[794] + l[843] + l[862] + l[869] + l[878] + l[888] + l[891] + l[908] + l[910] + l[929] + l[935] + l[940] + l[943] + l[946] + l[972] + l[981] + l[997] + l[1007] + l[1011] + l[1017] + l[1034] + l[1043] + l[1056] + l[1068] + l[1071] + l[1076] + l[1084] + l[1095] + l[1112] + l[1119] + l[1128] + l[1141] + l[1149] + l[1167] + l[1171] + l[1175] + l[1179] + l[1181] + l[1192] + l[1195] + l[1202] + l[1206] + l[1215] + l[1217] + l[1224] + l[1231] + l[1233] + l[1234] + l[1236] + l[1243] + l[1256] + l[1257] + l[1267] + l[1273] + l[1287] + l[1294] + l[1302] + l[1310] + l[1319] + l[1325] + l[1329] + l[1338] + l[1364] + l[1372] + l[1374] + l[1376]; // 0.03125
	assign val[7] = l[39] + l[43] + l[123] + l[158] + l[161] + l[164] + l[168] + l[174] + l[181] + l[225] + l[234] + l[238] + l[244] + l[253] + l[285] + l[298] + l[302] + l[318] + l[322] + l[341] + l[343] + l[357] + l[359] + l[364] + l[381] + l[383] + l[394] + l[406] + l[418] + l[423] + l[445] + l[467] + l[469] + l[476] + l[477] + l[482] + l[484] + l[485] + l[504] + l[513] + l[538] + l[542] + l[550] + l[558] + l[566] + l[571] + l[577] + l[596] + l[610] + l[614] + l[624] + l[651] + l[657] + l[661] + l[664] + l[667] + l[683] + l[689] + l[692] + l[696] + l[704] + l[707] + l[714] + l[719] + l[721] + l[722] + l[743] + l[745] + l[756] + l[759] + l[766] + l[768] + l[801] + l[818] + l[820] + l[830] + l[838] + l[841] + l[847] + l[851] + l[853] + l[873] + l[875] + l[886] + l[895] + l[897] + l[901] + l[905] + l[912] + l[918] + l[921] + l[924] + l[932] + l[934] + l[949] + l[955] + l[968] + l[971] + l[980] + l[984] + l[986] + l[990] + l[992] + l[995] + l[999] + l[1001] + l[1012] + l[1016] + l[1026] + l[1030] + l[1035] + l[1045] + l[1054] + l[1057] + l[1062] + l[1078] + l[1079] + l[1081] + l[1086] + l[1089] + l[1102] + l[1104] + l[1108] + l[1110] + l[1117] + l[1122] + l[1134] + l[1137] + l[1144] + l[1158] + l[1159] + l[1164] + l[1166] + l[1169] + l[1184] + l[1188] + l[1193] + l[1198] + l[1200] + l[1209] + l[1211] + l[1225] + l[1246] + l[1250] + l[1253] + l[1265] + l[1276] + l[1280] + l[1285] + l[1290] + l[1301] + l[1308] + l[1314] + l[1320] + l[1323] + l[1352] + l[1355] + l[1381] + l[1388] + l[1391] + l[1397] + l[1398]; // 0.0625
	assign val[8] = l[29] + l[30] + l[33] + l[51] + l[54] + l[63] + l[74] + l[81] + l[108] + l[127] + l[133] + l[135] + l[137] + l[145] + l[150] + l[162] + l[167] + l[187] + l[196] + l[199] + l[206] + l[211] + l[213] + l[220] + l[222] + l[230] + l[239] + l[241] + l[245] + l[255] + l[258] + l[260] + l[261] + l[267] + l[269] + l[277] + l[283] + l[286] + l[292] + l[295] + l[303] + l[305] + l[310] + l[323] + l[328] + l[330] + l[335] + l[338] + l[345] + l[346] + l[353] + l[361] + l[369] + l[377] + l[385] + l[393] + l[399] + l[410] + l[413] + l[415] + l[417] + l[426] + l[437] + l[455] + l[459] + l[472] + l[493] + l[496] + l[512] + l[516] + l[520] + l[524] + l[525] + l[532] + l[535] + l[539] + l[543] + l[546] + l[548] + l[552] + l[562] + l[563] + l[573] + l[581] + l[582] + l[591] + l[604] + l[619] + l[622] + l[626] + l[634] + l[643] + l[646] + l[658] + l[671] + l[674] + l[678] + l[694] + l[703] + l[711] + l[716] + l[731] + l[740] + l[754] + l[771] + l[773] + l[774] + l[781] + l[783] + l[786] + l[789] + l[797] + l[809] + l[813] + l[814] + l[817] + l[823] + l[825] + l[829] + l[835] + l[844] + l[854] + l[858] + l[860] + l[870] + l[880] + l[882] + l[885] + l[902] + l[911] + l[926] + l[928] + l[938] + l[939] + l[944] + l[950] + l[959] + l[960] + l[967] + l[1005] + l[1008] + l[1019] + l[1040] + l[1051] + l[1058] + l[1063] + l[1073] + l[1100] + l[1107] + l[1120] + l[1126] + l[1131] + l[1139] + l[1142] + l[1148] + l[1151] + l[1156] + l[1174] + l[1182] + l[1189] + l[1204] + l[1219] + l[1227] + l[1229] + l[1240] + l[1242] + l[1248] + l[1251] + l[1255] + l[1259] + l[1263] + l[1271] + l[1293] + l[1297] + l[1304] + l[1312] + l[1333] + l[1334] + l[1342] + l[1343] + l[1347] + l[1350] + l[1357] + l[1362] + l[1363] + l[1367] + l[1373] + l[1383] + l[1390]; // 0.125
	assign val[9] = l[6] + l[25] + l[40] + l[46] + l[58] + l[64] + l[66] + l[70] + l[73] + l[78] + l[83] + l[84] + l[90] + l[94] + l[97] + l[100] + l[102] + l[111] + l[115] + l[116] + l[120] + l[128] + l[130] + l[139] + l[142] + l[147] + l[148] + l[156] + l[163] + l[171] + l[177] + l[178] + l[182] + l[191] + l[193] + l[198] + l[208] + l[217] + l[223] + l[231] + l[251] + l[293] + l[319] + l[326] + l[334] + l[350] + l[367] + l[375] + l[380] + l[390] + l[396] + l[403] + l[428] + l[430] + l[435] + l[443] + l[454] + l[474] + l[478] + l[480] + l[488] + l[495] + l[503] + l[507] + l[556] + l[570] + l[595] + l[600] + l[618] + l[629] + l[632] + l[642] + l[648] + l[686] + l[724] + l[741] + l[744] + l[751] + l[776] + l[805] + l[808] + l[881] + l[920] + l[930] + l[964] + l[1031] + l[1038] + l[1042] + l[1065] + l[1114] + l[1123] + l[1214] + l[1324]; // 0.25
	assign val[10] = l[9] + l[17] + l[19] + l[22] + l[26] + l[31] + l[35] + l[36] + l[52] + l[88] + l[99] + l[401] + l[404] + l[434] + l[557] + l[583] + l[670]; // 0.5
	assign val[11] = l[2] + l[12] + l[42]; // 1.0
	assign val[12] = l[4] + l[8]; // 2.0
endmodule

module leaf_counter_6(input logic [0:1336] l, output logic [7:0] val [0:12]);
	assign val[0] = l[6] + l[12] + l[36] + l[48] + l[59] + l[63] + l[120] + l[125] + l[140] + l[147] + l[155] + l[163] + l[215] + l[267] + l[276] + l[281] + l[294] + l[297] + l[303] + l[312] + l[337] + l[339] + l[343] + l[363] + l[384] + l[392] + l[402] + l[410] + l[419] + l[432] + l[468] + l[476] + l[484] + l[492] + l[514] + l[517] + l[525] + l[559] + l[568] + l[583] + l[595] + l[600] + l[605] + l[627] + l[639] + l[661] + l[669] + l[683] + l[703] + l[717] + l[729] + l[732] + l[743] + l[777] + l[781] + l[807] + l[811] + l[821] + l[824] + l[835] + l[849] + l[854] + l[869] + l[874] + l[898] + l[948] + l[968] + l[977] + l[982] + l[1009] + l[1028] + l[1036] + l[1063] + l[1065] + l[1073] + l[1093] + l[1199] + l[1291] + l[1328]; // -0.25
	assign val[1] = l[0] + l[3] + l[10] + l[13] + l[14] + l[16] + l[22] + l[26] + l[28] + l[32] + l[41] + l[42] + l[44] + l[47] + l[51] + l[53] + l[56] + l[60] + l[62] + l[65] + l[68] + l[69] + l[73] + l[75] + l[78] + l[79] + l[82] + l[83] + l[86] + l[87] + l[93] + l[94] + l[97] + l[100] + l[102] + l[105] + l[108] + l[109] + l[115] + l[117] + l[124] + l[128] + l[130] + l[131] + l[136] + l[137] + l[142] + l[143] + l[145] + l[148] + l[149] + l[152] + l[154] + l[158] + l[161] + l[165] + l[167] + l[169] + l[171] + l[172] + l[174] + l[176] + l[179] + l[182] + l[184] + l[187] + l[192] + l[195] + l[196] + l[199] + l[200] + l[203] + l[207] + l[210] + l[211] + l[213] + l[218] + l[221] + l[223] + l[227] + l[229] + l[233] + l[234] + l[239] + l[241] + l[243] + l[244] + l[246] + l[247] + l[250] + l[257] + l[260] + l[263] + l[266] + l[268] + l[270] + l[271] + l[273] + l[283] + l[286] + l[287] + l[289] + l[296] + l[299] + l[302] + l[309] + l[314] + l[320] + l[321] + l[324] + l[327] + l[331] + l[336] + l[340] + l[345] + l[346] + l[348] + l[352] + l[357] + l[358] + l[360] + l[369] + l[370] + l[373] + l[378] + l[380] + l[386] + l[387] + l[393] + l[395] + l[396] + l[397] + l[405] + l[415] + l[418] + l[421] + l[423] + l[424] + l[431] + l[435] + l[440] + l[442] + l[444] + l[445] + l[448] + l[450] + l[451] + l[453] + l[461] + l[466] + l[470] + l[477] + l[482] + l[485] + l[488] + l[494] + l[496] + l[497] + l[500] + l[505] + l[506] + l[510] + l[516] + l[518] + l[519] + l[522] + l[527] + l[529] + l[532] + l[535] + l[538] + l[539] + l[541] + l[546] + l[550] + l[551] + l[557] + l[560] + l[561] + l[569] + l[572] + l[573] + l[575] + l[576] + l[578] + l[580] + l[582] + l[586] + l[592] + l[597] + l[604] + l[611] + l[612] + l[620] + l[624] + l[626] + l[629] + l[631] + l[632] + l[634] + l[637] + l[642] + l[646] + l[648] + l[656] + l[664] + l[668] + l[673] + l[674] + l[678] + l[679] + l[682] + l[685] + l[691] + l[694] + l[698] + l[706] + l[707] + l[711] + l[722] + l[724] + l[733] + l[736] + l[750] + l[752] + l[760] + l[762] + l[767] + l[768] + l[771] + l[774] + l[782] + l[793] + l[796] + l[797] + l[802] + l[804] + l[805] + l[808] + l[809] + l[813] + l[815] + l[820] + l[826] + l[829] + l[833] + l[838] + l[845] + l[851] + l[857] + l[861] + l[862] + l[867] + l[875] + l[876] + l[882] + l[885] + l[889] + l[890] + l[894] + l[903] + l[908] + l[912] + l[914] + l[918] + l[920] + l[924] + l[925] + l[928] + l[929] + l[930] + l[935] + l[938] + l[941] + l[944] + l[947] + l[950] + l[952] + l[960] + l[964] + l[969] + l[973] + l[980] + l[984] + l[986] + l[991] + l[993] + l[998] + l[1002] + l[1014] + l[1016] + l[1021] + l[1022] + l[1024] + l[1027] + l[1033] + l[1038] + l[1044] + l[1047] + l[1049] + l[1052] + l[1053] + l[1055] + l[1066] + l[1070] + l[1080] + l[1086] + l[1090] + l[1096] + l[1097] + l[1102] + l[1104] + l[1109] + l[1111] + l[1113] + l[1118] + l[1119] + l[1122] + l[1123] + l[1136] + l[1142] + l[1148] + l[1151] + l[1154] + l[1156] + l[1161] + l[1167] + l[1174] + l[1176] + l[1187] + l[1188] + l[1191] + l[1193] + l[1194] + l[1207] + l[1212] + l[1218] + l[1219] + l[1221] + l[1231] + l[1234] + l[1236] + l[1239] + l[1240] + l[1249] + l[1258] + l[1261] + l[1268] + l[1272] + l[1274] + l[1277] + l[1284] + l[1289] + l[1297] + l[1302] + l[1305] + l[1309] + l[1311] + l[1314] + l[1317] + l[1323] + l[1333]; // -0.125
	assign val[2] = l[19] + l[31] + l[34] + l[64] + l[116] + l[126] + l[133] + l[164] + l[188] + l[191] + l[193] + l[202] + l[212] + l[225] + l[249] + l[251] + l[254] + l[255] + l[258] + l[284] + l[305] + l[308] + l[311] + l[315] + l[334] + l[338] + l[341] + l[383] + l[388] + l[411] + l[414] + l[417] + l[429] + l[433] + l[456] + l[459] + l[464] + l[465] + l[472] + l[474] + l[490] + l[509] + l[530] + l[533] + l[542] + l[544] + l[555] + l[584] + l[590] + l[599] + l[606] + l[607] + l[616] + l[618] + l[622] + l[635] + l[651] + l[654] + l[658] + l[663] + l[666] + l[671] + l[677] + l[689] + l[704] + l[714] + l[727] + l[731] + l[737] + l[740] + l[745] + l[748] + l[754] + l[784] + l[791] + l[832] + l[836] + l[843] + l[844] + l[846] + l[855] + l[864] + l[865] + l[880] + l[897] + l[899] + l[915] + l[917] + l[923] + l[937] + l[958] + l[963] + l[972] + l[989] + l[997] + l[1001] + l[1003] + l[1005] + l[1026] + l[1030] + l[1035] + l[1041] + l[1057] + l[1061] + l[1064] + l[1074] + l[1076] + l[1081] + l[1105] + l[1110] + l[1128] + l[1131] + l[1134] + l[1140] + l[1145] + l[1152] + l[1158] + l[1164] + l[1165] + l[1172] + l[1183] + l[1200] + l[1204] + l[1205] + l[1220] + l[1223] + l[1226] + l[1232] + l[1246] + l[1253] + l[1255] + l[1265] + l[1271] + l[1280] + l[1292] + l[1294] + l[1296] + l[1308] + l[1316] + l[1322] + l[1326] + l[1329] + l[1332] + l[1334]; // -0.0625
	assign val[3] = l[58] + l[160] + l[280] + l[293] + l[304] + l[323] + l[350] + l[364] + l[377] + l[390] + l[401] + l[436] + l[441] + l[487] + l[588] + l[596] + l[602] + l[710] + l[751] + l[757] + l[778] + l[789] + l[799] + l[812] + l[818] + l[828] + l[841] + l[870] + l[878] + l[887] + l[922] + l[979] + l[994] + l[1011] + l[1040] + l[1046] + l[1062] + l[1072] + l[1082] + l[1092] + l[1094] + l[1116] + l[1120] + l[1126] + l[1179] + l[1181] + l[1197] + l[1202] + l[1209] + l[1229] + l[1245] + l[1278] + l[1285] + l[1287] + l[1299]; // -0.03125
	assign val[4] = l[80] + l[206] + l[230] + l[235] + l[238] + l[264] + l[328] + l[426] + l[469] + l[479] + l[493] + l[524] + l[623] + l[628] + l[645] + l[659] + l[680] + l[701] + l[715] + l[721] + l[758] + l[765] + l[776] + l[780] + l[783] + l[806] + l[852] + l[901] + l[910] + l[983] + l[1007] + l[1010] + l[1018] + l[1139] + l[1155] + l[1162] + l[1175] + l[1214] + l[1263] + l[1266] + l[1290] + l[1312] + l[1327]; // -0.015625
	assign val[5] = l[72] + l[111] + l[157] + l[275] + l[443] + l[481] + l[495] + l[501] + l[552] + l[577] + l[613] + l[614] + l[649] + l[693] + l[718] + l[755] + l[830] + l[871] + l[888] + l[893] + l[959] + l[967] + l[974] + l[981] + l[999] + l[1004] + l[1017] + l[1032] + l[1068] + l[1114] + l[1137] + l[1143] + l[1147] + l[1150] + l[1186] + l[1230] + l[1237] + l[1247] + l[1252] + l[1269] + l[1273] + l[1279] + l[1286] + l[1298] + l[1313] + l[1318] + l[1335]; // 0.015625
	assign val[6] = l[9] + l[156] + l[162] + l[197] + l[224] + l[269] + l[277] + l[298] + l[318] + l[329] + l[347] + l[354] + l[362] + l[400] + l[413] + l[420] + l[430] + l[437] + l[462] + l[502] + l[543] + l[547] + l[549] + l[571] + l[574] + l[587] + l[603] + l[621] + l[630] + l[647] + l[657] + l[672] + l[675] + l[686] + l[697] + l[699] + l[708] + l[712] + l[723] + l[744] + l[770] + l[795] + l[810] + l[816] + l[827] + l[834] + l[837] + l[847] + l[848] + l[860] + l[877] + l[904] + l[911] + l[939] + l[940] + l[942] + l[949] + l[951] + l[961] + l[965] + l[995] + l[1008] + l[1020] + l[1023] + l[1025] + l[1051] + l[1060] + l[1077] + l[1089] + l[1095] + l[1121] + l[1124] + l[1125] + l[1129] + l[1141] + l[1157] + l[1163] + l[1189] + l[1192] + l[1195] + l[1206] + l[1217] + l[1235] + l[1248] + l[1264] + l[1275] + l[1304] + l[1306] + l[1321] + l[1324] + l[1331]; // 0.03125
	assign val[7] = l[20] + l[25] + l[43] + l[55] + l[110] + l[144] + l[166] + l[177] + l[189] + l[216] + l[282] + l[300] + l[310] + l[316] + l[322] + l[335] + l[349] + l[359] + l[368] + l[372] + l[376] + l[394] + l[398] + l[409] + l[422] + l[438] + l[446] + l[455] + l[457] + l[467] + l[475] + l[478] + l[483] + l[486] + l[491] + l[498] + l[504] + l[508] + l[511] + l[523] + l[528] + l[534] + l[545] + l[558] + l[608] + l[617] + l[619] + l[638] + l[643] + l[644] + l[653] + l[681] + l[695] + l[716] + l[720] + l[730] + l[734] + l[738] + l[739] + l[741] + l[756] + l[763] + l[766] + l[775] + l[798] + l[800] + l[817] + l[819] + l[823] + l[839] + l[842] + l[859] + l[863] + l[868] + l[881] + l[891] + l[900] + l[906] + l[907] + l[916] + l[919] + l[934] + l[936] + l[946] + l[953] + l[956] + l[962] + l[978] + l[985] + l[987] + l[988] + l[990] + l[1000] + l[1006] + l[1013] + l[1037] + l[1042] + l[1050] + l[1058] + l[1067] + l[1075] + l[1091] + l[1100] + l[1103] + l[1112] + l[1117] + l[1130] + l[1135] + l[1144] + l[1153] + l[1173] + l[1182] + l[1215] + l[1224] + l[1227] + l[1228] + l[1238] + l[1241] + l[1242] + l[1257] + l[1267] + l[1270] + l[1288] + l[1295] + l[1307] + l[1310] + l[1325] + l[1330]; // 0.0625
	assign val[8] = l[5] + l[7] + l[37] + l[45] + l[66] + l[81] + l[84] + l[88] + l[101] + l[103] + l[129] + l[138] + l[141] + l[159] + l[178] + l[180] + l[185] + l[190] + l[208] + l[209] + l[214] + l[219] + l[228] + l[232] + l[240] + l[245] + l[248] + l[253] + l[256] + l[261] + l[279] + l[285] + l[290] + l[295] + l[306] + l[313] + l[317] + l[319] + l[332] + l[344] + l[361] + l[375] + l[382] + l[389] + l[391] + l[399] + l[412] + l[427] + l[428] + l[434] + l[447] + l[449] + l[460] + l[463] + l[473] + l[480] + l[489] + l[507] + l[513] + l[526] + l[537] + l[553] + l[556] + l[566] + l[570] + l[579] + l[585] + l[594] + l[598] + l[601] + l[609] + l[625] + l[636] + l[650] + l[662] + l[665] + l[667] + l[670] + l[676] + l[684] + l[687] + l[690] + l[692] + l[696] + l[700] + l[702] + l[709] + l[728] + l[747] + l[749] + l[759] + l[764] + l[779] + l[785] + l[787] + l[790] + l[792] + l[801] + l[803] + l[814] + l[825] + l[831] + l[840] + l[853] + l[866] + l[872] + l[879] + l[886] + l[892] + l[902] + l[909] + l[921] + l[927] + l[933] + l[955] + l[966] + l[971] + l[992] + l[996] + l[1031] + l[1039] + l[1045] + l[1048] + l[1059] + l[1069] + l[1078] + l[1083] + l[1088] + l[1106] + l[1115] + l[1132] + l[1138] + l[1146] + l[1149] + l[1160] + l[1166] + l[1169] + l[1178] + l[1180] + l[1185] + l[1196] + l[1201] + l[1203] + l[1210] + l[1213] + l[1222] + l[1233] + l[1244] + l[1251] + l[1256] + l[1262] + l[1276] + l[1282] + l[1283] + l[1293] + l[1300] + l[1303] + l[1315] + l[1319] + l[1336]; // 0.125
	assign val[9] = l[21] + l[23] + l[27] + l[29] + l[35] + l[39] + l[40] + l[49] + l[52] + l[54] + l[57] + l[67] + l[71] + l[74] + l[76] + l[85] + l[89] + l[96] + l[98] + l[113] + l[127] + l[132] + l[134] + l[135] + l[139] + l[150] + l[151] + l[170] + l[173] + l[175] + l[183] + l[186] + l[194] + l[198] + l[205] + l[217] + l[226] + l[242] + l[252] + l[272] + l[274] + l[278] + l[292] + l[301] + l[307] + l[326] + l[333] + l[342] + l[351] + l[355] + l[356] + l[365] + l[367] + l[381] + l[385] + l[404] + l[408] + l[416] + l[454] + l[458] + l[471] + l[499] + l[503] + l[520] + l[531] + l[548] + l[563] + l[589] + l[615] + l[640] + l[652] + l[655] + l[660] + l[719] + l[726] + l[773] + l[786] + l[896] + l[943] + l[975] + l[1012] + l[1019] + l[1034] + l[1085] + l[1101] + l[1108] + l[1127] + l[1171] + l[1198] + l[1259]; // 0.25
	assign val[10] = l[11] + l[15] + l[17] + l[18] + l[24] + l[33] + l[46] + l[50] + l[61] + l[70] + l[77] + l[92] + l[104] + l[106] + l[107] + l[112] + l[122] + l[153] + l[168] + l[201] + l[231] + l[236] + l[330] + l[439] + l[554]; // 0.5
	assign val[11] = l[1] + l[30] + l[38] + l[90] + l[91] + l[119]; // 1.0
	assign val[12] = l[2] + l[4] + l[8]; // 2.0
endmodule

module leaf_counter_7(input logic [0:1279] l, output logic [7:0] val [0:12]);
	assign val[0] = l[12] + l[21] + l[24] + l[30] + l[37] + l[50] + l[54] + l[56] + l[69] + l[73] + l[84] + l[87] + l[88] + l[92] + l[94] + l[99] + l[101] + l[111] + l[120] + l[146] + l[155] + l[156] + l[162] + l[175] + l[178] + l[185] + l[186] + l[203] + l[207] + l[218] + l[222] + l[240] + l[247] + l[265] + l[270] + l[275] + l[277] + l[282] + l[288] + l[300] + l[315] + l[320] + l[328] + l[342] + l[344] + l[346] + l[364] + l[368] + l[378] + l[380] + l[386] + l[388] + l[399] + l[405] + l[408] + l[410] + l[412] + l[417] + l[420] + l[426] + l[441] + l[445] + l[453] + l[455] + l[458] + l[475] + l[478] + l[489] + l[492] + l[501] + l[505] + l[510] + l[517] + l[520] + l[531] + l[540] + l[551] + l[558] + l[560] + l[561] + l[573] + l[583] + l[592] + l[604] + l[623] + l[628] + l[638] + l[639] + l[660] + l[666] + l[676] + l[689] + l[691] + l[697] + l[719] + l[726] + l[731] + l[749] + l[764] + l[789] + l[793] + l[799] + l[820] + l[824] + l[841] + l[846] + l[853] + l[855] + l[875] + l[908] + l[917] + l[925] + l[936] + l[940] + l[961] + l[965] + l[980] + l[983] + l[998] + l[1006] + l[1009] + l[1011] + l[1015] + l[1022] + l[1024] + l[1028] + l[1064] + l[1077] + l[1094] + l[1117] + l[1127] + l[1133] + l[1139] + l[1161] + l[1166] + l[1180] + l[1206] + l[1214] + l[1218] + l[1219] + l[1224] + l[1257] + l[1278]; // -0.25
	assign val[1] = l[0] + l[3] + l[10] + l[17] + l[18] + l[20] + l[23] + l[25] + l[26] + l[28] + l[33] + l[34] + l[36] + l[38] + l[40] + l[42] + l[44] + l[47] + l[49] + l[55] + l[58] + l[60] + l[63] + l[65] + l[67] + l[68] + l[71] + l[72] + l[74] + l[76] + l[81] + l[85] + l[89] + l[90] + l[95] + l[97] + l[102] + l[104] + l[112] + l[115] + l[116] + l[117] + l[118] + l[121] + l[124] + l[125] + l[129] + l[130] + l[133] + l[136] + l[140] + l[142] + l[145] + l[147] + l[150] + l[154] + l[158] + l[161] + l[164] + l[166] + l[169] + l[171] + l[172] + l[174] + l[183] + l[187] + l[188] + l[191] + l[192] + l[194] + l[196] + l[198] + l[210] + l[212] + l[214] + l[216] + l[219] + l[229] + l[232] + l[244] + l[249] + l[252] + l[254] + l[255] + l[259] + l[264] + l[268] + l[273] + l[276] + l[280] + l[291] + l[302] + l[303] + l[305] + l[307] + l[311] + l[312] + l[319] + l[331] + l[333] + l[336] + l[339] + l[354] + l[357] + l[359] + l[361] + l[363] + l[367] + l[372] + l[376] + l[379] + l[384] + l[389] + l[391] + l[395] + l[396] + l[403] + l[419] + l[421] + l[424] + l[431] + l[435] + l[437] + l[443] + l[449] + l[456] + l[459] + l[461] + l[466] + l[469] + l[481] + l[483] + l[484] + l[490] + l[494] + l[498] + l[500] + l[509] + l[514] + l[516] + l[519] + l[528] + l[529] + l[533] + l[535] + l[538] + l[544] + l[546] + l[549] + l[566] + l[572] + l[577] + l[579] + l[581] + l[587] + l[589] + l[596] + l[599] + l[603] + l[609] + l[611] + l[618] + l[624] + l[626] + l[634] + l[642] + l[651] + l[657] + l[664] + l[668] + l[675] + l[681] + l[692] + l[693] + l[696] + l[700] + l[702] + l[705] + l[712] + l[718] + l[720] + l[724] + l[729] + l[730] + l[737] + l[739] + l[743] + l[747] + l[748] + l[755] + l[760] + l[762] + l[763] + l[767] + l[770] + l[771] + l[776] + l[777] + l[778] + l[783] + l[798] + l[805] + l[807] + l[809] + l[810] + l[812] + l[814] + l[817] + l[822] + l[829] + l[833] + l[836] + l[839] + l[845] + l[847] + l[850] + l[852] + l[860] + l[861] + l[862] + l[866] + l[873] + l[878] + l[880] + l[888] + l[891] + l[896] + l[904] + l[911] + l[913] + l[919] + l[927] + l[929] + l[933] + l[938] + l[939] + l[942] + l[947] + l[952] + l[960] + l[962] + l[964] + l[972] + l[974] + l[977] + l[979] + l[984] + l[990] + l[999] + l[1019] + l[1030] + l[1033] + l[1040] + l[1042] + l[1045] + l[1046] + l[1050] + l[1055] + l[1056] + l[1062] + l[1073] + l[1080] + l[1086] + l[1091] + l[1101] + l[1104] + l[1108] + l[1112] + l[1113] + l[1122] + l[1123] + l[1126] + l[1130] + l[1132] + l[1154] + l[1156] + l[1163] + l[1169] + l[1189] + l[1197] + l[1198] + l[1200] + l[1204] + l[1212] + l[1217] + l[1225] + l[1236] + l[1243] + l[1245] + l[1253] + l[1262] + l[1263] + l[1267] + l[1275]; // -0.125
	assign val[2] = l[5] + l[6] + l[13] + l[31] + l[83] + l[109] + l[110] + l[122] + l[126] + l[143] + l[148] + l[152] + l[159] + l[163] + l[176] + l[181] + l[197] + l[199] + l[225] + l[236] + l[237] + l[242] + l[245] + l[257] + l[267] + l[281] + l[284] + l[287] + l[294] + l[298] + l[299] + l[321] + l[343] + l[347] + l[350] + l[352] + l[355] + l[369] + l[387] + l[397] + l[400] + l[411] + l[413] + l[429] + l[434] + l[464] + l[474] + l[485] + l[487] + l[502] + l[511] + l[536] + l[541] + l[552] + l[562] + l[568] + l[569] + l[576] + l[578] + l[600] + l[614] + l[629] + l[646] + l[648] + l[650] + l[671] + l[686] + l[687] + l[690] + l[709] + l[714] + l[723] + l[727] + l[734] + l[751] + l[753] + l[769] + l[779] + l[795] + l[800] + l[815] + l[823] + l[842] + l[856] + l[857] + l[868] + l[879] + l[885] + l[892] + l[895] + l[903] + l[918] + l[922] + l[935] + l[944] + l[945] + l[951] + l[955] + l[970] + l[976] + l[988] + l[991] + l[1001] + l[1013] + l[1018] + l[1034] + l[1053] + l[1058] + l[1065] + l[1067] + l[1072] + l[1076] + l[1082] + l[1085] + l[1088] + l[1098] + l[1103] + l[1116] + l[1128] + l[1134] + l[1138] + l[1140] + l[1153] + l[1165] + l[1171] + l[1174] + l[1178] + l[1179] + l[1182] + l[1183] + l[1186] + l[1190] + l[1193] + l[1203] + l[1207] + l[1209] + l[1221] + l[1227] + l[1233] + l[1240] + l[1255] + l[1261] + l[1277]; // -0.0625
	assign val[3] = l[139] + l[157] + l[189] + l[250] + l[261] + l[296] + l[317] + l[322] + l[324] + l[365] + l[383] + l[401] + l[404] + l[416] + l[427] + l[438] + l[450] + l[472] + l[504] + l[521] + l[548] + l[555] + l[556] + l[598] + l[607] + l[610] + l[619] + l[632] + l[640] + l[653] + l[656] + l[658] + l[667] + l[677] + l[679] + l[699] + l[708] + l[711] + l[721] + l[738] + l[745] + l[772] + l[774] + l[782] + l[784] + l[788] + l[790] + l[792] + l[797] + l[819] + l[827] + l[844] + l[870] + l[882] + l[890] + l[900] + l[916] + l[948] + l[956] + l[959] + l[967] + l[981] + l[993] + l[1010] + l[1037] + l[1039] + l[1051] + l[1074] + l[1099] + l[1110] + l[1136] + l[1147] + l[1173] + l[1215] + l[1232] + l[1239] + l[1247] + l[1259] + l[1271] + l[1273] + l[1276]; // -0.03125
	assign val[4] = l[53] + l[100] + l[107] + l[123] + l[184] + l[211] + l[239] + l[266] + l[285] + l[304] + l[335] + l[393] + l[406] + l[414] + l[496] + l[506] + l[513] + l[525] + l[526] + l[582] + l[612] + l[636] + l[643] + l[716] + l[811] + l[831] + l[854] + l[932] + l[950] + l[986] + l[992] + l[1000] + l[1007] + l[1025] + l[1043] + l[1057] + l[1069] + l[1105] + l[1155] + l[1188] + l[1194] + l[1230] + l[1249] + l[1252] + l[1269]; // -0.015625
	assign val[5] = l[103] + l[173] + l[224] + l[306] + l[314] + l[345] + l[432] + l[465] + l[468] + l[503] + l[534] + l[554] + l[563] + l[565] + l[591] + l[605] + l[659] + l[662] + l[674] + l[715] + l[746] + l[804] + l[806] + l[864] + l[886] + l[897] + l[920] + l[957] + l[968] + l[989] + l[1031] + l[1041] + l[1047] + l[1049] + l[1060] + l[1083] + l[1111] + l[1160] + l[1162] + l[1213] + l[1216] + l[1241] + l[1254]; // 0.015625
	assign val[6] = l[15] + l[51] + l[61] + l[78] + l[80] + l[86] + l[131] + l[153] + l[165] + l[168] + l[179] + l[182] + l[215] + l[258] + l[283] + l[292] + l[308] + l[318] + l[327] + l[366] + l[373] + l[382] + l[394] + l[407] + l[409] + l[418] + l[423] + l[436] + l[446] + l[471] + l[497] + l[512] + l[527] + l[542] + l[543] + l[570] + l[575] + l[584] + l[586] + l[588] + l[620] + l[649] + l[654] + l[661] + l[665] + l[670] + l[722] + l[736] + l[744] + l[750] + l[766] + l[773] + l[775] + l[813] + l[834] + l[837] + l[872] + l[889] + l[894] + l[898] + l[907] + l[915] + l[931] + l[934] + l[943] + l[946] + l[958] + l[973] + l[982] + l[1016] + l[1020] + l[1026] + l[1029] + l[1044] + l[1052] + l[1063] + l[1081] + l[1087] + l[1096] + l[1106] + l[1121] + l[1125] + l[1129] + l[1131] + l[1137] + l[1149] + l[1164] + l[1211] + l[1231] + l[1238] + l[1258] + l[1270]; // 0.03125
	assign val[7] = l[39] + l[48] + l[66] + l[113] + l[190] + l[195] + l[200] + l[201] + l[204] + l[220] + l[226] + l[230] + l[243] + l[248] + l[256] + l[274] + l[301] + l[313] + l[323] + l[332] + l[337] + l[351] + l[360] + l[362] + l[425] + l[430] + l[440] + l[444] + l[454] + l[488] + l[499] + l[507] + l[515] + l[532] + l[537] + l[547] + l[567] + l[571] + l[597] + l[602] + l[615] + l[617] + l[625] + l[627] + l[635] + l[644] + l[669] + l[684] + l[703] + l[710] + l[728] + l[741] + l[796] + l[803] + l[821] + l[826] + l[828] + l[830] + l[840] + l[843] + l[851] + l[858] + l[869] + l[877] + l[881] + l[901] + l[910] + l[912] + l[926] + l[963] + l[975] + l[978] + l[987] + l[1004] + l[1032] + l[1038] + l[1054] + l[1059] + l[1068] + l[1079] + l[1093] + l[1097] + l[1100] + l[1109] + l[1119] + l[1120] + l[1141] + l[1145] + l[1152] + l[1158] + l[1181] + l[1184] + l[1187] + l[1191] + l[1199] + l[1226] + l[1242] + l[1248] + l[1251] + l[1256] + l[1264] + l[1272] + l[1274] + l[1279]; // 0.0625
	assign val[8] = l[35] + l[62] + l[77] + l[91] + l[96] + l[98] + l[132] + l[138] + l[151] + l[170] + l[180] + l[202] + l[205] + l[213] + l[228] + l[241] + l[253] + l[262] + l[263] + l[272] + l[278] + l[279] + l[286] + l[297] + l[310] + l[316] + l[325] + l[330] + l[334] + l[338] + l[341] + l[349] + l[358] + l[370] + l[381] + l[392] + l[402] + l[415] + l[428] + l[433] + l[448] + l[451] + l[452] + l[457] + l[467] + l[470] + l[473] + l[477] + l[480] + l[495] + l[518] + l[522] + l[524] + l[545] + l[553] + l[557] + l[559] + l[580] + l[593] + l[595] + l[601] + l[606] + l[608] + l[613] + l[622] + l[631] + l[637] + l[645] + l[647] + l[655] + l[663] + l[673] + l[678] + l[682] + l[685] + l[688] + l[694] + l[695] + l[698] + l[701] + l[706] + l[707] + l[713] + l[754] + l[756] + l[780] + l[781] + l[785] + l[787] + l[791] + l[808] + l[816] + l[818] + l[832] + l[838] + l[848] + l[863] + l[871] + l[874] + l[883] + l[887] + l[893] + l[902] + l[905] + l[906] + l[914] + l[924] + l[928] + l[930] + l[937] + l[954] + l[969] + l[994] + l[996] + l[1008] + l[1017] + l[1035] + l[1061] + l[1070] + l[1071] + l[1084] + l[1115] + l[1135] + l[1142] + l[1150] + l[1167] + l[1172] + l[1177] + l[1185] + l[1192] + l[1195] + l[1201] + l[1202] + l[1205] + l[1208] + l[1222] + l[1228] + l[1235] + l[1250]; // 0.125
	assign val[9] = l[22] + l[32] + l[41] + l[46] + l[52] + l[64] + l[70] + l[75] + l[82] + l[93] + l[106] + l[108] + l[114] + l[134] + l[141] + l[149] + l[160] + l[167] + l[193] + l[206] + l[209] + l[217] + l[221] + l[223] + l[231] + l[233] + l[235] + l[238] + l[246] + l[260] + l[269] + l[289] + l[293] + l[295] + l[326] + l[353] + l[375] + l[422] + l[447] + l[463] + l[486] + l[491] + l[508] + l[523] + l[564] + l[574] + l[585] + l[590] + l[630] + l[680] + l[704] + l[732] + l[740] + l[759] + l[849] + l[865] + l[884] + l[899] + l[921] + l[941] + l[949] + l[971] + l[1002] + l[1036] + l[1048] + l[1089] + l[1118] + l[1124] + l[1146] + l[1176] + l[1229] + l[1237] + l[1244] + l[1265]; // 0.25
	assign val[10] = l[1] + l[9] + l[16] + l[19] + l[27] + l[29] + l[43] + l[59] + l[79] + l[119] + l[127] + l[128] + l[137] + l[144] + l[177] + l[234] + l[309] + l[356] + l[717] + l[742] + l[757]; // 0.5
	assign val[11] = l[2] + l[7] + l[11] + l[14] + l[105]; // 1.0
	assign val[12] = l[4] + l[8]; // 2.0
endmodule

module leaf_counter_8(input logic [0:1497] l, output logic [7:0] val [0:12]);
	assign val[0] = l[2] + l[48] + l[64] + l[96] + l[140] + l[167] + l[172] + l[206] + l[294] + l[366] + l[412] + l[429] + l[593] + l[597] + l[639] + l[665] + l[668] + l[690] + l[727] + l[733] + l[782] + l[793] + l[811] + l[822] + l[841] + l[855] + l[1077] + l[1345] + l[1385] + l[1426] + l[1437]; // -0.25
	assign val[1] = l[0] + l[1] + l[4] + l[8] + l[16] + l[18] + l[22] + l[24] + l[32] + l[33] + l[34] + l[36] + l[40] + l[42] + l[44] + l[49] + l[50] + l[54] + l[56] + l[65] + l[66] + l[68] + l[72] + l[80] + l[82] + l[86] + l[88] + l[97] + l[99] + l[101] + l[104] + l[110] + l[112] + l[117] + l[120] + l[126] + l[132] + l[136] + l[141] + l[143] + l[144] + l[150] + l[152] + l[160] + l[168] + l[173] + l[174] + l[176] + l[188] + l[191] + l[192] + l[199] + l[204] + l[217] + l[222] + l[227] + l[232] + l[236] + l[252] + l[254] + l[258] + l[260] + l[263] + l[266] + l[268] + l[277] + l[280] + l[284] + l[287] + l[288] + l[292] + l[295] + l[300] + l[316] + l[323] + l[327] + l[331] + l[333] + l[335] + l[351] + l[356] + l[358] + l[359] + l[377] + l[378] + l[382] + l[385] + l[386] + l[402] + l[404] + l[406] + l[417] + l[422] + l[426] + l[428] + l[438] + l[444] + l[445] + l[452] + l[459] + l[461] + l[466] + l[469] + l[475] + l[478] + l[483] + l[485] + l[497] + l[499] + l[505] + l[507] + l[517] + l[519] + l[523] + l[533] + l[538] + l[540] + l[541] + l[544] + l[552] + l[560] + l[570] + l[572] + l[580] + l[587] + l[591] + l[596] + l[600] + l[609] + l[614] + l[628] + l[631] + l[638] + l[646] + l[648] + l[653] + l[659] + l[670] + l[677] + l[681] + l[689] + l[703] + l[706] + l[707] + l[720] + l[722] + l[730] + l[731] + l[736] + l[737] + l[761] + l[774] + l[777] + l[780] + l[786] + l[787] + l[789] + l[795] + l[796] + l[799] + l[800] + l[805] + l[809] + l[819] + l[824] + l[835] + l[840] + l[852] + l[861] + l[864] + l[872] + l[885] + l[886] + l[889] + l[892] + l[896] + l[903] + l[908] + l[916] + l[920] + l[924] + l[936] + l[946] + l[970] + l[972] + l[974] + l[976] + l[977] + l[979] + l[984] + l[995] + l[1003] + l[1027] + l[1029] + l[1032] + l[1040] + l[1045] + l[1046] + l[1070] + l[1080] + l[1082] + l[1091] + l[1102] + l[1107] + l[1125] + l[1126] + l[1140] + l[1146] + l[1151] + l[1158] + l[1172] + l[1191] + l[1193] + l[1202] + l[1212] + l[1215] + l[1234] + l[1244] + l[1253] + l[1258] + l[1264] + l[1275] + l[1276] + l[1278] + l[1282] + l[1299] + l[1300] + l[1304] + l[1306] + l[1310] + l[1314] + l[1318] + l[1322] + l[1334] + l[1346] + l[1349] + l[1352] + l[1364] + l[1372] + l[1373] + l[1393] + l[1408] + l[1411] + l[1416] + l[1439] + l[1443] + l[1451] + l[1453] + l[1475] + l[1479] + l[1481] + l[1487] + l[1491]; // -0.125
	assign val[2] = l[13] + l[26] + l[52] + l[59] + l[62] + l[76] + l[85] + l[91] + l[94] + l[128] + l[134] + l[166] + l[178] + l[184] + l[195] + l[196] + l[208] + l[212] + l[216] + l[224] + l[230] + l[238] + l[240] + l[242] + l[248] + l[265] + l[275] + l[290] + l[298] + l[304] + l[313] + l[322] + l[329] + l[341] + l[343] + l[347] + l[367] + l[373] + l[390] + l[396] + l[399] + l[403] + l[409] + l[418] + l[424] + l[430] + l[432] + l[436] + l[468] + l[501] + l[506] + l[515] + l[525] + l[537] + l[547] + l[555] + l[557] + l[581] + l[582] + l[601] + l[611] + l[621] + l[629] + l[632] + l[640] + l[641] + l[649] + l[656] + l[671] + l[674] + l[688] + l[693] + l[696] + l[699] + l[715] + l[728] + l[734] + l[743] + l[748] + l[752] + l[755] + l[757] + l[768] + l[781] + l[784] + l[801] + l[815] + l[823] + l[827] + l[842] + l[843] + l[850] + l[856] + l[857] + l[873] + l[879] + l[890] + l[898] + l[912] + l[927] + l[929] + l[940] + l[953] + l[955] + l[959] + l[962] + l[980] + l[990] + l[992] + l[1002] + l[1008] + l[1015] + l[1020] + l[1022] + l[1026] + l[1035] + l[1043] + l[1049] + l[1050] + l[1053] + l[1057] + l[1060] + l[1062] + l[1065] + l[1069] + l[1073] + l[1078] + l[1090] + l[1098] + l[1109] + l[1111] + l[1116] + l[1121] + l[1123] + l[1133] + l[1135] + l[1143] + l[1153] + l[1163] + l[1164] + l[1169] + l[1174] + l[1179] + l[1189] + l[1198] + l[1219] + l[1221] + l[1232] + l[1240] + l[1242] + l[1250] + l[1254] + l[1260] + l[1262] + l[1266] + l[1281] + l[1284] + l[1288] + l[1291] + l[1303] + l[1324] + l[1326] + l[1331] + l[1333] + l[1335] + l[1337] + l[1340] + l[1360] + l[1367] + l[1374] + l[1375] + l[1378] + l[1383] + l[1388] + l[1396] + l[1402] + l[1405] + l[1419] + l[1423] + l[1430] + l[1436] + l[1447] + l[1448] + l[1460] + l[1468] + l[1469] + l[1473] + l[1495] + l[1497]; // -0.0625
	assign val[3] = l[17] + l[69] + l[71] + l[102] + l[130] + l[149] + l[154] + l[171] + l[177] + l[219] + l[235] + l[247] + l[256] + l[259] + l[278] + l[296] + l[307] + l[350] + l[353] + l[375] + l[389] + l[440] + l[458] + l[488] + l[493] + l[510] + l[530] + l[564] + l[565] + l[573] + l[575] + l[577] + l[579] + l[586] + l[604] + l[607] + l[610] + l[617] + l[634] + l[661] + l[666] + l[679] + l[683] + l[692] + l[712] + l[713] + l[724] + l[740] + l[745] + l[753] + l[770] + l[775] + l[804] + l[806] + l[833] + l[837] + l[882] + l[893] + l[901] + l[905] + l[931] + l[933] + l[935] + l[947] + l[965] + l[985] + l[987] + l[997] + l[1011] + l[1017] + l[1038] + l[1089] + l[1092] + l[1095] + l[1104] + l[1114] + l[1129] + l[1130] + l[1145] + l[1155] + l[1156] + l[1170] + l[1194] + l[1206] + l[1209] + l[1225] + l[1228] + l[1237] + l[1272] + l[1277] + l[1283] + l[1312] + l[1317] + l[1319] + l[1351] + l[1354] + l[1371] + l[1384] + l[1387] + l[1399] + l[1421] + l[1425] + l[1428] + l[1438] + l[1452] + l[1455] + l[1465] + l[1476] + l[1480] + l[1484]; // -0.03125
	assign val[4] = l[20] + l[28] + l[39] + l[74] + l[100] + l[145] + l[180] + l[251] + l[283] + l[395] + l[407] + l[411] + l[414] + l[447] + l[453] + l[465] + l[471] + l[481] + l[492] + l[528] + l[542] + l[549] + l[636] + l[642] + l[657] + l[709] + l[719] + l[773] + l[812] + l[846] + l[854] + l[880] + l[938] + l[943] + l[956] + l[957] + l[999] + l[1013] + l[1031] + l[1047] + l[1058] + l[1101] + l[1106] + l[1127] + l[1160] + l[1173] + l[1177] + l[1201] + l[1217] + l[1226] + l[1247] + l[1294] + l[1301] + l[1358] + l[1365] + l[1369] + l[1381] + l[1424] + l[1450] + l[1459] + l[1462] + l[1485] + l[1488]; // -0.015625
	assign val[5] = l[207] + l[225] + l[274] + l[352] + l[379] + l[398] + l[401] + l[439] + l[451] + l[464] + l[509] + l[526] + l[558] + l[563] + l[618] + l[622] + l[633] + l[652] + l[660] + l[723] + l[741] + l[766] + l[769] + l[778] + l[792] + l[825] + l[844] + l[911] + l[921] + l[941] + l[952] + l[981] + l[1001] + l[1005] + l[1023] + l[1067] + l[1079] + l[1085] + l[1087] + l[1099] + l[1175] + l[1181] + l[1185] + l[1203] + l[1210] + l[1222] + l[1231] + l[1235] + l[1257] + l[1259] + l[1271] + l[1297] + l[1305] + l[1327] + l[1347] + l[1368] + l[1382] + l[1442] + l[1444] + l[1467] + l[1477] + l[1482] + l[1486] + l[1489]; // 0.015625
	assign val[6] = l[67] + l[73] + l[113] + l[114] + l[137] + l[146] + l[151] + l[205] + l[220] + l[233] + l[237] + l[249] + l[255] + l[269] + l[293] + l[301] + l[321] + l[328] + l[337] + l[339] + l[342] + l[365] + l[392] + l[421] + l[460] + l[470] + l[512] + l[521] + l[531] + l[534] + l[543] + l[559] + l[561] + l[574] + l[590] + l[613] + l[695] + l[697] + l[701] + l[721] + l[738] + l[746] + l[758] + l[767] + l[816] + l[828] + l[836] + l[847] + l[849] + l[851] + l[860] + l[871] + l[874] + l[883] + l[888] + l[917] + l[925] + l[934] + l[937] + l[949] + l[961] + l[969] + l[973] + l[1025] + l[1036] + l[1061] + l[1075] + l[1094] + l[1097] + l[1103] + l[1118] + l[1120] + l[1124] + l[1134] + l[1148] + l[1150] + l[1165] + l[1168] + l[1176] + l[1178] + l[1195] + l[1218] + l[1224] + l[1233] + l[1236] + l[1238] + l[1243] + l[1273] + l[1274] + l[1338] + l[1342] + l[1380] + l[1398] + l[1407] + l[1413] + l[1415] + l[1422] + l[1431] + l[1433] + l[1435] + l[1466] + l[1470] + l[1474] + l[1492]; // 0.03125
	assign val[7] = l[23] + l[37] + l[51] + l[87] + l[93] + l[105] + l[107] + l[108] + l[111] + l[116] + l[119] + l[133] + l[179] + l[182] + l[185] + l[190] + l[214] + l[228] + l[231] + l[246] + l[264] + l[267] + l[289] + l[297] + l[306] + l[320] + l[344] + l[354] + l[384] + l[387] + l[391] + l[397] + l[405] + l[413] + l[416] + l[427] + l[431] + l[433] + l[437] + l[456] + l[462] + l[474] + l[476] + l[484] + l[502] + l[508] + l[524] + l[527] + l[535] + l[548] + l[551] + l[576] + l[602] + l[606] + l[608] + l[630] + l[637] + l[647] + l[654] + l[662] + l[669] + l[676] + l[682] + l[685] + l[687] + l[694] + l[700] + l[708] + l[710] + l[716] + l[718] + l[744] + l[747] + l[750] + l[754] + l[756] + l[759] + l[762] + l[772] + l[779] + l[790] + l[797] + l[803] + l[807] + l[821] + l[832] + l[834] + l[839] + l[862] + l[884] + l[891] + l[900] + l[902] + l[907] + l[909] + l[913] + l[914] + l[926] + l[930] + l[939] + l[944] + l[948] + l[954] + l[960] + l[966] + l[967] + l[988] + l[989] + l[993] + l[996] + l[1000] + l[1016] + l[1018] + l[1021] + l[1037] + l[1041] + l[1044] + l[1051] + l[1054] + l[1063] + l[1064] + l[1068] + l[1083] + l[1088] + l[1100] + l[1108] + l[1128] + l[1136] + l[1141] + l[1144] + l[1147] + l[1157] + l[1161] + l[1171] + l[1188] + l[1199] + l[1207] + l[1220] + l[1227] + l[1249] + l[1252] + l[1255] + l[1267] + l[1279] + l[1280] + l[1285] + l[1287] + l[1290] + l[1292] + l[1295] + l[1302] + l[1307] + l[1321] + l[1328] + l[1332] + l[1336] + l[1339] + l[1353] + l[1357] + l[1359] + l[1361] + l[1363] + l[1370] + l[1376] + l[1379] + l[1389] + l[1391] + l[1401] + l[1404] + l[1420] + l[1427] + l[1429] + l[1456] + l[1461] + l[1464] + l[1471] + l[1478] + l[1483] + l[1493] + l[1496]; // 0.0625
	assign val[8] = l[5] + l[6] + l[9] + l[25] + l[35] + l[41] + l[57] + l[60] + l[78] + l[83] + l[84] + l[89] + l[95] + l[121] + l[125] + l[127] + l[129] + l[135] + l[139] + l[153] + l[155] + l[157] + l[159] + l[161] + l[163] + l[165] + l[169] + l[170] + l[181] + l[187] + l[193] + l[194] + l[197] + l[200] + l[203] + l[209] + l[210] + l[223] + l[234] + l[239] + l[241] + l[243] + l[244] + l[257] + l[261] + l[271] + l[273] + l[279] + l[282] + l[285] + l[291] + l[299] + l[311] + l[318] + l[325] + l[334] + l[345] + l[348] + l[349] + l[355] + l[357] + l[360] + l[368] + l[369] + l[372] + l[374] + l[380] + l[388] + l[408] + l[415] + l[419] + l[425] + l[434] + l[442] + l[450] + l[454] + l[463] + l[472] + l[479] + l[482] + l[486] + l[487] + l[491] + l[494] + l[495] + l[500] + l[513] + l[516] + l[529] + l[532] + l[546] + l[554] + l[556] + l[566] + l[567] + l[569] + l[571] + l[578] + l[588] + l[589] + l[595] + l[599] + l[603] + l[605] + l[612] + l[620] + l[626] + l[627] + l[635] + l[650] + l[651] + l[655] + l[658] + l[663] + l[667] + l[672] + l[673] + l[678] + l[680] + l[684] + l[686] + l[704] + l[705] + l[711] + l[717] + l[732] + l[735] + l[739] + l[742] + l[751] + l[764] + l[776] + l[783] + l[788] + l[791] + l[808] + l[818] + l[826] + l[829] + l[845] + l[848] + l[853] + l[858] + l[865] + l[866] + l[870] + l[875] + l[878] + l[895] + l[904] + l[910] + l[918] + l[923] + l[932] + l[942] + l[950] + l[951] + l[958] + l[963] + l[978] + l[982] + l[986] + l[998] + l[1006] + l[1014] + l[1019] + l[1024] + l[1030] + l[1034] + l[1039] + l[1048] + l[1052] + l[1055] + l[1056] + l[1059] + l[1066] + l[1071] + l[1072] + l[1074] + l[1076] + l[1081] + l[1084] + l[1086] + l[1093] + l[1096] + l[1105] + l[1113] + l[1115] + l[1117] + l[1119] + l[1131] + l[1132] + l[1137] + l[1138] + l[1154] + l[1162] + l[1167] + l[1180] + l[1183] + l[1186] + l[1197] + l[1200] + l[1208] + l[1211] + l[1216] + l[1223] + l[1230] + l[1239] + l[1246] + l[1248] + l[1256] + l[1261] + l[1263] + l[1268] + l[1270] + l[1289] + l[1296] + l[1311] + l[1315] + l[1320] + l[1323] + l[1330] + l[1341] + l[1344] + l[1350] + l[1366] + l[1377] + l[1386] + l[1395] + l[1406] + l[1410] + l[1414] + l[1417] + l[1432] + l[1434] + l[1440] + l[1446] + l[1449] + l[1457] + l[1490] + l[1494]; // 0.125
	assign val[9] = l[10] + l[14] + l[19] + l[30] + l[45] + l[47] + l[53] + l[58] + l[63] + l[70] + l[75] + l[77] + l[79] + l[90] + l[92] + l[103] + l[106] + l[109] + l[118] + l[123] + l[124] + l[131] + l[142] + l[147] + l[148] + l[156] + l[164] + l[175] + l[183] + l[186] + l[189] + l[198] + l[201] + l[213] + l[215] + l[218] + l[226] + l[229] + l[245] + l[250] + l[276] + l[281] + l[286] + l[303] + l[310] + l[312] + l[314] + l[324] + l[326] + l[330] + l[338] + l[340] + l[346] + l[361] + l[363] + l[371] + l[376] + l[393] + l[394] + l[400] + l[410] + l[420] + l[435] + l[441] + l[443] + l[448] + l[455] + l[457] + l[467] + l[473] + l[490] + l[503] + l[511] + l[522] + l[536] + l[539] + l[550] + l[553] + l[562] + l[568] + l[583] + l[615] + l[623] + l[643] + l[675] + l[691] + l[698] + l[702] + l[714] + l[726] + l[729] + l[749] + l[765] + l[798] + l[810] + l[813] + l[831] + l[838] + l[863] + l[867] + l[881] + l[906] + l[968] + l[994] + l[1010] + l[1012] + l[1042] + l[1149] + l[1205] + l[1293] + l[1308] + l[1325] + l[1355] + l[1356] + l[1390] + l[1463]; // 0.25
	assign val[10] = l[3] + l[12] + l[27] + l[29] + l[31] + l[38] + l[43] + l[46] + l[55] + l[61] + l[115] + l[138] + l[221] + l[309] + l[364] + l[514] + l[584] + l[644]; // 0.5
	assign val[11] = l[7] + l[11] + l[15] + l[21]; // 1.0
	assign val[12] = 0; // 2.0
endmodule

module leaf_counter_9(input logic [0:1347] l, output logic [7:0] val [0:12]);
	assign val[0] = l[24] + l[28] + l[53] + l[81] + l[93] + l[110] + l[119] + l[123] + l[129] + l[133] + l[145] + l[155] + l[159] + l[171] + l[173] + l[196] + l[207] + l[210] + l[223] + l[234] + l[237] + l[240] + l[245] + l[250] + l[260] + l[266] + l[275] + l[277] + l[296] + l[305] + l[308] + l[319] + l[321] + l[325] + l[341] + l[351] + l[352] + l[357] + l[367] + l[368] + l[377] + l[394] + l[421] + l[426] + l[429] + l[442] + l[468] + l[477] + l[492] + l[496] + l[507] + l[519] + l[531] + l[535] + l[558] + l[563] + l[572] + l[591] + l[602] + l[608] + l[612] + l[617] + l[623] + l[626] + l[636] + l[644] + l[655] + l[661] + l[669] + l[676] + l[687] + l[697] + l[700] + l[718] + l[725] + l[748] + l[754] + l[761] + l[820] + l[828] + l[846] + l[869] + l[885] + l[909] + l[948] + l[982] + l[1041] + l[1052] + l[1104] + l[1111] + l[1182] + l[1292]; // -0.25
	assign val[1] = l[0] + l[8] + l[16] + l[20] + l[25] + l[27] + l[30] + l[34] + l[38] + l[41] + l[45] + l[49] + l[57] + l[60] + l[64] + l[68] + l[70] + l[72] + l[80] + l[83] + l[87] + l[89] + l[98] + l[99] + l[109] + l[111] + l[112] + l[114] + l[115] + l[117] + l[122] + l[125] + l[130] + l[132] + l[136] + l[137] + l[141] + l[143] + l[148] + l[152] + l[161] + l[164] + l[165] + l[174] + l[176] + l[177] + l[179] + l[180] + l[182] + l[184] + l[187] + l[188] + l[191] + l[194] + l[198] + l[201] + l[205] + l[206] + l[208] + l[211] + l[213] + l[215] + l[218] + l[221] + l[224] + l[226] + l[229] + l[232] + l[243] + l[244] + l[246] + l[251] + l[252] + l[254] + l[256] + l[263] + l[279] + l[280] + l[282] + l[283] + l[287] + l[292] + l[295] + l[297] + l[300] + l[302] + l[303] + l[306] + l[310] + l[312] + l[315] + l[323] + l[327] + l[329] + l[336] + l[345] + l[354] + l[356] + l[358] + l[363] + l[365] + l[371] + l[373] + l[379] + l[382] + l[384] + l[385] + l[391] + l[396] + l[397] + l[400] + l[402] + l[403] + l[409] + l[412] + l[417] + l[419] + l[424] + l[427] + l[431] + l[433] + l[436] + l[440] + l[448] + l[450] + l[454] + l[459] + l[460] + l[461] + l[463] + l[466] + l[478] + l[484] + l[490] + l[501] + l[510] + l[513] + l[515] + l[517] + l[524] + l[526] + l[532] + l[539] + l[541] + l[548] + l[554] + l[556] + l[565] + l[566] + l[574] + l[580] + l[584] + l[588] + l[590] + l[614] + l[629] + l[634] + l[651] + l[674] + l[680] + l[683] + l[686] + l[690] + l[693] + l[703] + l[707] + l[708] + l[710] + l[714] + l[717] + l[729] + l[732] + l[736] + l[738] + l[742] + l[755] + l[757] + l[768] + l[775] + l[780] + l[787] + l[791] + l[795] + l[797] + l[798] + l[802] + l[804] + l[811] + l[812] + l[817] + l[818] + l[821] + l[825] + l[826] + l[832] + l[839] + l[840] + l[849] + l[853] + l[859] + l[870] + l[873] + l[886] + l[891] + l[898] + l[900] + l[906] + l[908] + l[910] + l[914] + l[919] + l[921] + l[929] + l[937] + l[947] + l[951] + l[953] + l[954] + l[961] + l[965] + l[969] + l[971] + l[978] + l[980] + l[981] + l[992] + l[994] + l[997] + l[1003] + l[1005] + l[1009] + l[1020] + l[1027] + l[1035] + l[1037] + l[1049] + l[1053] + l[1058] + l[1059] + l[1063] + l[1069] + l[1071] + l[1075] + l[1081] + l[1085] + l[1088] + l[1094] + l[1106] + l[1115] + l[1117] + l[1123] + l[1128] + l[1132] + l[1136] + l[1139] + l[1143] + l[1148] + l[1150] + l[1154] + l[1165] + l[1168] + l[1172] + l[1185] + l[1186] + l[1187] + l[1193] + l[1198] + l[1201] + l[1204] + l[1205] + l[1215] + l[1221] + l[1229] + l[1230] + l[1236] + l[1241] + l[1255] + l[1260] + l[1265] + l[1273] + l[1274] + l[1279] + l[1280] + l[1286] + l[1287] + l[1289] + l[1293] + l[1300] + l[1302] + l[1314] + l[1317] + l[1323] + l[1325] + l[1328] + l[1333] + l[1343] + l[1344]; // -0.125
	assign val[2] = l[4] + l[47] + l[52] + l[55] + l[76] + l[79] + l[91] + l[94] + l[95] + l[100] + l[101] + l[103] + l[106] + l[134] + l[149] + l[151] + l[154] + l[166] + l[172] + l[175] + l[178] + l[212] + l[238] + l[239] + l[253] + l[257] + l[281] + l[284] + l[309] + l[320] + l[322] + l[326] + l[330] + l[332] + l[335] + l[350] + l[353] + l[366] + l[375] + l[389] + l[393] + l[414] + l[434] + l[456] + l[469] + l[470] + l[472] + l[476] + l[487] + l[494] + l[495] + l[500] + l[504] + l[505] + l[525] + l[527] + l[534] + l[537] + l[553] + l[559] + l[561] + l[570] + l[573] + l[582] + l[585] + l[587] + l[592] + l[596] + l[601] + l[605] + l[619] + l[621] + l[631] + l[666] + l[677] + l[691] + l[699] + l[701] + l[719] + l[724] + l[733] + l[760] + l[763] + l[765] + l[769] + l[785] + l[805] + l[806] + l[823] + l[836] + l[841] + l[842] + l[854] + l[862] + l[865] + l[876] + l[915] + l[917] + l[923] + l[925] + l[933] + l[938] + l[941] + l[943] + l[945] + l[957] + l[959] + l[976] + l[984] + l[990] + l[998] + l[1007] + l[1008] + l[1014] + l[1043] + l[1045] + l[1066] + l[1090] + l[1093] + l[1096] + l[1126] + l[1141] + l[1144] + l[1153] + l[1170] + l[1174] + l[1176] + l[1188] + l[1191] + l[1218] + l[1220] + l[1224] + l[1227] + l[1239] + l[1243] + l[1247] + l[1257] + l[1259] + l[1262] + l[1268] + l[1278] + l[1281] + l[1284] + l[1290] + l[1294] + l[1311] + l[1318] + l[1320] + l[1330] + l[1339]; // -0.0625
	assign val[3] = l[2] + l[46] + l[75] + l[127] + l[147] + l[216] + l[233] + l[247] + l[313] + l[333] + l[337] + l[360] + l[362] + l[438] + l[441] + l[480] + l[483] + l[516] + l[522] + l[544] + l[562] + l[577] + l[594] + l[613] + l[627] + l[637] + l[641] + l[654] + l[660] + l[670] + l[722] + l[726] + l[728] + l[731] + l[741] + l[788] + l[831] + l[833] + l[856] + l[880] + l[884] + l[889] + l[972] + l[989] + l[996] + l[1001] + l[1013] + l[1017] + l[1023] + l[1029] + l[1033] + l[1047] + l[1067] + l[1074] + l[1079] + l[1084] + l[1100] + l[1102] + l[1105] + l[1108] + l[1116] + l[1137] + l[1160] + l[1171] + l[1195] + l[1210] + l[1211] + l[1238] + l[1242] + l[1276] + l[1297] + l[1307] + l[1312] + l[1316] + l[1322] + l[1329] + l[1332] + l[1334] + l[1340]; // -0.03125
	assign val[4] = l[17] + l[29] + l[113] + l[156] + l[168] + l[195] + l[220] + l[274] + l[290] + l[369] + l[388] + l[458] + l[497] + l[555] + l[609] + l[610] + l[622] + l[625] + l[635] + l[640] + l[667] + l[682] + l[698] + l[713] + l[744] + l[782] + l[875] + l[883] + l[894] + l[896] + l[928] + l[963] + l[983] + l[1042] + l[1060] + l[1076] + l[1083] + l[1109] + l[1112] + l[1114] + l[1124] + l[1129] + l[1135] + l[1146] + l[1177] + l[1184] + l[1214] + l[1234] + l[1246] + l[1253] + l[1270] + l[1272] + l[1298] + l[1336] + l[1342] + l[1347]; // -0.015625
	assign val[5] = l[37] + l[204] + l[241] + l[271] + l[346] + l[372] + l[395] + l[432] + l[449] + l[464] + l[506] + l[560] + l[564] + l[578] + l[581] + l[600] + l[606] + l[638] + l[656] + l[684] + l[706] + l[709] + l[716] + l[745] + l[762] + l[781] + l[786] + l[807] + l[827] + l[837] + l[838] + l[895] + l[926] + l[930] + l[964] + l[966] + l[968] + l[1018] + l[1080] + l[1120] + l[1147] + l[1163] + l[1189] + l[1226] + l[1231] + l[1235] + l[1258] + l[1269] + l[1275] + l[1309] + l[1327]; // 0.015625
	assign val[6] = l[21] + l[31] + l[54] + l[82] + l[126] + l[138] + l[200] + l[214] + l[222] + l[242] + l[286] + l[301] + l[328] + l[364] + l[411] + l[423] + l[428] + l[437] + l[453] + l[485] + l[489] + l[503] + l[508] + l[521] + l[528] + l[533] + l[549] + l[567] + l[576] + l[589] + l[616] + l[618] + l[649] + l[657] + l[668] + l[689] + l[715] + l[721] + l[735] + l[740] + l[743] + l[750] + l[752] + l[773] + l[799] + l[810] + l[824] + l[852] + l[857] + l[858] + l[871] + l[872] + l[881] + l[882] + l[887] + l[897] + l[903] + l[905] + l[912] + l[942] + l[946] + l[950] + l[958] + l[973] + l[1006] + l[1012] + l[1015] + l[1016] + l[1024] + l[1031] + l[1072] + l[1082] + l[1089] + l[1103] + l[1107] + l[1122] + l[1164] + l[1173] + l[1175] + l[1181] + l[1190] + l[1192] + l[1194] + l[1199] + l[1206] + l[1212] + l[1216] + l[1219] + l[1222] + l[1223] + l[1245] + l[1251] + l[1283] + l[1299] + l[1313] + l[1321] + l[1331] + l[1335]; // 0.03125
	assign val[7] = l[13] + l[14] + l[50] + l[58] + l[62] + l[67] + l[85] + l[88] + l[92] + l[104] + l[135] + l[146] + l[153] + l[158] + l[181] + l[185] + l[186] + l[189] + l[190] + l[217] + l[219] + l[231] + l[235] + l[255] + l[278] + l[293] + l[316] + l[318] + l[324] + l[349] + l[355] + l[378] + l[381] + l[383] + l[390] + l[399] + l[401] + l[406] + l[408] + l[415] + l[420] + l[457] + l[465] + l[467] + l[473] + l[479] + l[502] + l[536] + l[550] + l[552] + l[583] + l[597] + l[599] + l[607] + l[620] + l[643] + l[663] + l[671] + l[678] + l[685] + l[694] + l[705] + l[712] + l[723] + l[730] + l[759] + l[766] + l[770] + l[772] + l[800] + l[813] + l[829] + l[835] + l[848] + l[851] + l[855] + l[861] + l[874] + l[902] + l[907] + l[918] + l[920] + l[927] + l[932] + l[935] + l[944] + l[952] + l[956] + l[960] + l[975] + l[977] + l[987] + l[1004] + l[1021] + l[1025] + l[1034] + l[1038] + l[1040] + l[1044] + l[1046] + l[1048] + l[1056] + l[1068] + l[1073] + l[1078] + l[1092] + l[1099] + l[1101] + l[1110] + l[1118] + l[1125] + l[1127] + l[1131] + l[1138] + l[1140] + l[1145] + l[1151] + l[1152] + l[1155] + l[1158] + l[1166] + l[1169] + l[1179] + l[1202] + l[1203] + l[1208] + l[1209] + l[1217] + l[1232] + l[1240] + l[1264] + l[1267] + l[1271] + l[1282] + l[1285] + l[1301] + l[1310] + l[1319] + l[1345] + l[1346]; // 0.0625
	assign val[8] = l[6] + l[9] + l[10] + l[22] + l[35] + l[44] + l[61] + l[78] + l[84] + l[96] + l[108] + l[118] + l[121] + l[124] + l[131] + l[139] + l[160] + l[162] + l[170] + l[183] + l[193] + l[203] + l[209] + l[259] + l[261] + l[264] + l[267] + l[269] + l[272] + l[276] + l[289] + l[291] + l[307] + l[311] + l[334] + l[339] + l[342] + l[361] + l[370] + l[376] + l[386] + l[387] + l[398] + l[404] + l[410] + l[418] + l[439] + l[443] + l[444] + l[447] + l[451] + l[471] + l[474] + l[481] + l[482] + l[486] + l[491] + l[493] + l[499] + l[509] + l[518] + l[520] + l[530] + l[538] + l[540] + l[546] + l[557] + l[569] + l[571] + l[575] + l[579] + l[586] + l[593] + l[595] + l[611] + l[615] + l[624] + l[632] + l[639] + l[648] + l[652] + l[673] + l[675] + l[681] + l[696] + l[702] + l[711] + l[734] + l[746] + l[774] + l[778] + l[783] + l[789] + l[792] + l[794] + l[809] + l[815] + l[822] + l[830] + l[845] + l[863] + l[867] + l[868] + l[877] + l[888] + l[892] + l[899] + l[916] + l[931] + l[939] + l[962] + l[967] + l[985] + l[995] + l[999] + l[1000] + l[1010] + l[1019] + l[1032] + l[1054] + l[1061] + l[1065] + l[1077] + l[1086] + l[1091] + l[1097] + l[1113] + l[1119] + l[1134] + l[1156] + l[1162] + l[1178] + l[1197] + l[1200] + l[1213] + l[1225] + l[1228] + l[1237] + l[1248] + l[1254] + l[1261] + l[1288] + l[1295] + l[1296] + l[1304] + l[1326] + l[1338] + l[1341]; // 0.125
	assign val[9] = l[18] + l[32] + l[36] + l[40] + l[48] + l[51] + l[65] + l[66] + l[71] + l[77] + l[90] + l[97] + l[102] + l[107] + l[128] + l[142] + l[144] + l[150] + l[157] + l[163] + l[192] + l[197] + l[199] + l[225] + l[227] + l[228] + l[236] + l[249] + l[262] + l[265] + l[273] + l[285] + l[299] + l[314] + l[331] + l[338] + l[343] + l[347] + l[359] + l[374] + l[405] + l[416] + l[435] + l[446] + l[462] + l[488] + l[512] + l[529] + l[543] + l[545] + l[568] + l[642] + l[646] + l[647] + l[650] + l[659] + l[664] + l[672] + l[692] + l[727] + l[739] + l[749] + l[764] + l[801] + l[814] + l[843] + l[860] + l[878] + l[890] + l[893] + l[901] + l[904] + l[913] + l[924] + l[934] + l[986] + l[991] + l[1022] + l[1026] + l[1030] + l[1064] + l[1157] + l[1180] + l[1196] + l[1207] + l[1249] + l[1252] + l[1263] + l[1308] + l[1337]; // 0.25
	assign val[10] = l[1] + l[5] + l[23] + l[42] + l[56] + l[63] + l[73] + l[74] + l[86] + l[105] + l[116] + l[167] + l[268] + l[407] + l[498] + l[658] + l[790] + l[844]; // 0.5
	assign val[11] = l[3] + l[7] + l[11] + l[15] + l[19] + l[33] + l[43] + l[59]; // 1.0
	assign val[12] = l[12]; // 2.0
endmodule